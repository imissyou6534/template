module accel_control(
  input         clock,
  input         reset,
  input         io_ap_done,
  input         io_pool_finish_edge,
  output        io_conv_finish,
  output [31:0] io_reg0,
  output [31:0] io_reg1,
  output [31:0] io_reg2,
  output [31:0] io_reg3,
  output [31:0] io_reg4,
  output [31:0] io_reg5,
  output [31:0] io_reg6,
  output [31:0] io_reg7,
  output [31:0] io_reg8,
  output [31:0] io_reg9,
  output [31:0] io_reg10,
  output        io_yolo_finish,
  output        io_resize_load
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
`endif // RANDOMIZE_REG_INIT
  reg  yolo_finish; // @[control.scala 40:28]
  reg  io_yolo_finish_REG; // @[utils.scala 10:17]
  reg  ap_done_up_REG; // @[utils.scala 10:17]
  wire  ap_done_up = ~ap_done_up_REG & io_ap_done; // @[utils.scala 10:27]
  reg [3:0] c2f_cnt; // @[control.scala 46:26]
  wire  _c2f_shortcut_T = c2f_cnt == 4'h1; // @[control.scala 49:52]
  wire  _c2f_shortcut_T_1 = c2f_cnt == 4'h2; // @[control.scala 49:76]
  wire  _c2f_shortcut_T_2 = c2f_cnt == 4'h3; // @[control.scala 49:100]
  wire  _c2f_shortcut_T_3 = c2f_cnt == 4'h0; // @[control.scala 49:124]
  wire  _c2f_shortcut_T_6 = c2f_cnt == 4'h7; // @[control.scala 49:198]
  wire  c2f_shortcut = _c2f_shortcut_T | (_c2f_shortcut_T_1 | (_c2f_shortcut_T_2 | _c2f_shortcut_T_3)); // @[Mux.scala 101:16]
  reg [4:0] current_layer; // @[control.scala 52:32]
  wire  cur_layer_sel_0 = current_layer == 5'h0; // @[control.scala 58:81]
  wire  cur_layer_sel_1 = current_layer == 5'h1; // @[control.scala 58:81]
  wire  cur_layer_sel_2 = current_layer == 5'h2; // @[control.scala 58:81]
  wire  cur_layer_sel_3 = current_layer == 5'h3; // @[control.scala 58:81]
  wire  cur_layer_sel_4 = current_layer == 5'h4; // @[control.scala 58:81]
  wire  cur_layer_sel_5 = current_layer == 5'h5; // @[control.scala 58:81]
  wire  cur_layer_sel_6 = current_layer == 5'h6; // @[control.scala 58:81]
  wire  cur_layer_sel_7 = current_layer == 5'h7; // @[control.scala 58:81]
  wire  cur_layer_sel_8 = current_layer == 5'h8; // @[control.scala 58:81]
  wire  cur_layer_sel_9 = current_layer == 5'h9; // @[control.scala 58:81]
  wire  cur_layer_sel_10 = current_layer == 5'ha; // @[control.scala 58:81]
  wire  cur_layer_sel_11 = current_layer == 5'hb; // @[control.scala 58:81]
  wire  cur_layer_sel_12 = current_layer == 5'hc; // @[control.scala 58:81]
  wire  cur_layer_sel_13 = current_layer == 5'hd; // @[control.scala 58:81]
  wire  cur_layer_sel_14 = current_layer == 5'he; // @[control.scala 58:81]
  wire  cur_layer_sel_15 = current_layer == 5'hf; // @[control.scala 58:81]
  wire  cur_layer_sel_16 = current_layer == 5'h10; // @[control.scala 58:81]
  wire  cur_layer_sel_17 = current_layer == 5'h11; // @[control.scala 58:81]
  wire  cur_layer_sel_18 = current_layer == 5'h12; // @[control.scala 58:81]
  wire  cur_layer_sel_19 = current_layer == 5'h13; // @[control.scala 58:81]
  wire  cur_layer_sel_20 = current_layer == 5'h14; // @[control.scala 58:81]
  wire  cur_layer_sel_21 = current_layer == 5'h15; // @[control.scala 58:81]
  wire [6:0] _current_layer_cout_T = cur_layer_sel_21 ? 7'h50 : 7'h0; // @[Mux.scala 101:16]
  wire [6:0] _current_layer_cout_T_1 = cur_layer_sel_20 ? 7'h50 : _current_layer_cout_T; // @[Mux.scala 101:16]
  wire [6:0] _current_layer_cout_T_2 = cur_layer_sel_19 ? 7'h50 : _current_layer_cout_T_1; // @[Mux.scala 101:16]
  wire [6:0] _current_layer_cout_T_3 = cur_layer_sel_18 ? 7'h40 : _current_layer_cout_T_2; // @[Mux.scala 101:16]
  wire [6:0] _current_layer_cout_T_4 = cur_layer_sel_17 ? 7'h40 : _current_layer_cout_T_3; // @[Mux.scala 101:16]
  wire [6:0] _current_layer_cout_T_5 = cur_layer_sel_16 ? 7'h40 : _current_layer_cout_T_4; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_6 = cur_layer_sel_15 ? 9'h100 : {{2'd0}, _current_layer_cout_T_5}; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_7 = cur_layer_sel_14 ? 9'h80 : _current_layer_cout_T_6; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_8 = cur_layer_sel_13 ? 9'h80 : _current_layer_cout_T_7; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_9 = cur_layer_sel_12 ? 9'h40 : _current_layer_cout_T_8; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_10 = cur_layer_sel_11 ? 9'h40 : _current_layer_cout_T_9; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_11 = cur_layer_sel_10 ? 9'h80 : _current_layer_cout_T_10; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_12 = cur_layer_sel_9 ? 9'h100 : _current_layer_cout_T_11; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_13 = cur_layer_sel_8 ? 9'h100 : _current_layer_cout_T_12; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_14 = cur_layer_sel_7 ? 9'h100 : _current_layer_cout_T_13; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_15 = cur_layer_sel_6 ? 9'h80 : _current_layer_cout_T_14; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_16 = cur_layer_sel_5 ? 9'h80 : _current_layer_cout_T_15; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_17 = cur_layer_sel_4 ? 9'h40 : _current_layer_cout_T_16; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_18 = cur_layer_sel_3 ? 9'h40 : _current_layer_cout_T_17; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_19 = cur_layer_sel_2 ? 9'h20 : _current_layer_cout_T_18; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_20 = cur_layer_sel_1 ? 9'h20 : _current_layer_cout_T_19; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cout_T_21 = cur_layer_sel_0 ? 9'h10 : _current_layer_cout_T_20; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T = cur_layer_sel_21 ? 9'h100 : 9'h0; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_1 = cur_layer_sel_20 ? 9'h80 : _current_layer_cin_T; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_2 = cur_layer_sel_19 ? 9'h40 : _current_layer_cin_T_1; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_3 = cur_layer_sel_18 ? 9'h100 : _current_layer_cin_T_2; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_4 = cur_layer_sel_17 ? 9'h80 : _current_layer_cin_T_3; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_5 = cur_layer_sel_16 ? 9'h40 : _current_layer_cin_T_4; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_6 = cur_layer_sel_15 ? 9'h180 : _current_layer_cin_T_5; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_7 = cur_layer_sel_14 ? 9'h80 : _current_layer_cin_T_6; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_8 = cur_layer_sel_13 ? 9'hc0 : _current_layer_cin_T_7; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_9 = cur_layer_sel_12 ? 9'h40 : _current_layer_cin_T_8; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_10 = cur_layer_sel_11 ? 9'hc0 : _current_layer_cin_T_9; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_11 = cur_layer_sel_10 ? 9'h180 : _current_layer_cin_T_10; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_12 = cur_layer_sel_9 ? 9'h100 : _current_layer_cin_T_11; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_13 = cur_layer_sel_8 ? 9'h100 : _current_layer_cin_T_12; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_14 = cur_layer_sel_7 ? 9'h80 : _current_layer_cin_T_13; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_15 = cur_layer_sel_6 ? 9'h80 : _current_layer_cin_T_14; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_16 = cur_layer_sel_5 ? 9'h40 : _current_layer_cin_T_15; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_17 = cur_layer_sel_4 ? 9'h40 : _current_layer_cin_T_16; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_18 = cur_layer_sel_3 ? 9'h20 : _current_layer_cin_T_17; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_19 = cur_layer_sel_2 ? 9'h20 : _current_layer_cin_T_18; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_20 = cur_layer_sel_1 ? 9'h10 : _current_layer_cin_T_19; // @[Mux.scala 101:16]
  wire [8:0] _current_layer_cin_T_21 = cur_layer_sel_0 ? 9'h8 : _current_layer_cin_T_20; // @[Mux.scala 101:16]
  wire  _current_layer_repeats_T_1 = cur_layer_sel_20 | cur_layer_sel_21; // @[Mux.scala 101:16]
  wire  _current_layer_repeats_T_14 = cur_layer_sel_7 | (cur_layer_sel_8 | (cur_layer_sel_9 | (cur_layer_sel_10 | (
    cur_layer_sel_11 | (cur_layer_sel_12 | (cur_layer_sel_13 | (cur_layer_sel_14 | (cur_layer_sel_15 | (cur_layer_sel_16
     | (cur_layer_sel_17 | (cur_layer_sel_18 | (cur_layer_sel_19 | (cur_layer_sel_20 | cur_layer_sel_21))))))))))))); // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_15 = cur_layer_sel_6 ? 2'h2 : {{1'd0}, _current_layer_repeats_T_14}; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_16 = cur_layer_sel_5 ? 2'h1 : _current_layer_repeats_T_15; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_17 = cur_layer_sel_4 ? 2'h2 : _current_layer_repeats_T_16; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_18 = cur_layer_sel_3 ? 2'h1 : _current_layer_repeats_T_17; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_19 = cur_layer_sel_2 ? 2'h1 : _current_layer_repeats_T_18; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_20 = cur_layer_sel_1 ? 2'h1 : _current_layer_repeats_T_19; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_repeats_T_21 = cur_layer_sel_0 ? 2'h1 : _current_layer_repeats_T_20; // @[Mux.scala 101:16]
  wire  _current_layer_sel_T_9 = cur_layer_sel_12 | cur_layer_sel_13; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_10 = cur_layer_sel_11 ? 2'h2 : {{1'd0}, _current_layer_sel_T_9}; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_11 = cur_layer_sel_10 ? 2'h1 : _current_layer_sel_T_10; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_12 = cur_layer_sel_9 ? 2'h0 : _current_layer_sel_T_11; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_13 = cur_layer_sel_8 ? 2'h0 : _current_layer_sel_T_12; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_14 = cur_layer_sel_7 ? 2'h0 : _current_layer_sel_T_13; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_15 = cur_layer_sel_6 ? 2'h1 : _current_layer_sel_T_14; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_16 = cur_layer_sel_5 ? 2'h1 : _current_layer_sel_T_15; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_17 = cur_layer_sel_4 ? 2'h2 : _current_layer_sel_T_16; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_18 = cur_layer_sel_3 ? 2'h2 : _current_layer_sel_T_17; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_19 = cur_layer_sel_2 ? 2'h3 : _current_layer_sel_T_18; // @[Mux.scala 101:16]
  wire [1:0] _current_layer_sel_T_20 = cur_layer_sel_1 ? 2'h3 : _current_layer_sel_T_19; // @[Mux.scala 101:16]
  wire [2:0] current_layer_sel = cur_layer_sel_0 ? 3'h4 : {{1'd0}, _current_layer_sel_T_20}; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T = cur_layer_sel_21 ? 3'h4 : 3'h0; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_1 = cur_layer_sel_20 ? 3'h4 : _current_model_code_T; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_2 = cur_layer_sel_19 ? 3'h4 : _current_model_code_T_1; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_3 = cur_layer_sel_18 ? 3'h3 : _current_model_code_T_2; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_4 = cur_layer_sel_17 ? 3'h3 : _current_model_code_T_3; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_5 = cur_layer_sel_16 ? 3'h3 : _current_model_code_T_4; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_6 = cur_layer_sel_15 ? 3'h1 : _current_model_code_T_5; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_7 = cur_layer_sel_14 ? 3'h0 : _current_model_code_T_6; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_8 = cur_layer_sel_13 ? 3'h1 : _current_model_code_T_7; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_9 = cur_layer_sel_12 ? 3'h0 : _current_model_code_T_8; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_10 = cur_layer_sel_11 ? 3'h1 : _current_model_code_T_9; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_11 = cur_layer_sel_10 ? 3'h1 : _current_model_code_T_10; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_12 = cur_layer_sel_9 ? 3'h2 : _current_model_code_T_11; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_13 = cur_layer_sel_8 ? 3'h1 : _current_model_code_T_12; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_14 = cur_layer_sel_7 ? 3'h0 : _current_model_code_T_13; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_15 = cur_layer_sel_6 ? 3'h1 : _current_model_code_T_14; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_16 = cur_layer_sel_5 ? 3'h0 : _current_model_code_T_15; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_17 = cur_layer_sel_4 ? 3'h1 : _current_model_code_T_16; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_18 = cur_layer_sel_3 ? 3'h0 : _current_model_code_T_17; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_19 = cur_layer_sel_2 ? 3'h1 : _current_model_code_T_18; // @[Mux.scala 101:16]
  wire [2:0] _current_model_code_T_20 = cur_layer_sel_1 ? 3'h0 : _current_model_code_T_19; // @[Mux.scala 101:16]
  wire [2:0] current_model_code = cur_layer_sel_0 ? 3'h0 : _current_model_code_T_20; // @[Mux.scala 101:16]
  reg  conv_finish; // @[control.scala 71:30]
  wire  current_layer_is_conv = current_model_code == 3'h0; // @[control.scala 75:52]
  wire  current_layer_is_c2f = current_model_code == 3'h1; // @[control.scala 76:51]
  wire  current_layer_is_sppf = current_model_code == 3'h2; // @[control.scala 77:52]
  wire  current_layer_is_detect_box = current_model_code == 3'h3; // @[control.scala 78:58]
  wire  current_layer_is_detect_cls = current_model_code == 3'h4; // @[control.scala 79:58]
  reg [4:0] current_layer_next; // @[control.scala 81:37]
  reg  current_layer_is_c2f_next; // @[control.scala 83:44]
  wire  _c2f_cnt_T = current_layer != current_layer_next; // @[control.scala 85:35]
  wire [3:0] _c2f_cnt_T_4 = c2f_cnt + 4'h1; // @[control.scala 85:135]
  wire [2:0] current_layer_repeats = {{1'd0}, _current_layer_repeats_T_21}; // @[control.scala 55:37 66:27]
  wire [5:0] _conv_number_in_c2f_T = {current_layer_repeats, 3'h0}; // @[control.scala 88:49]
  reg [4:0] conv_cnt_in_c2f; // @[control.scala 90:34]
  wire [4:0] conv_number_in_c2f = _conv_number_in_c2f_T[4:0]; // @[control.scala 86:34 88:24]
  wire [4:0] _conv_cnt_in_c2f_T_2 = conv_number_in_c2f - 5'h1; // @[control.scala 91:108]
  wire  _conv_cnt_in_c2f_T_3 = conv_cnt_in_c2f == _conv_cnt_in_c2f_T_2; // @[control.scala 91:84]
  wire [4:0] _conv_cnt_in_c2f_T_5 = conv_cnt_in_c2f + 5'h1; // @[control.scala 91:137]
  reg [2:0] cnt_in_sppf; // @[control.scala 93:30]
  wire  _cnt_in_sppf_T_1 = cnt_in_sppf == 3'h1; // @[control.scala 94:77]
  wire [2:0] _cnt_in_sppf_T_3 = cnt_in_sppf + 3'h1; // @[control.scala 94:118]
  reg [2:0] cnt_in_detect_box; // @[control.scala 96:36]
  wire  _cnt_in_detect_box_T_1 = cnt_in_detect_box == 3'h2; // @[control.scala 97:95]
  wire [2:0] _cnt_in_detect_box_T_3 = cnt_in_detect_box + 3'h1; // @[control.scala 97:148]
  reg [2:0] cnt_in_detect_cls; // @[control.scala 99:36]
  wire  _cnt_in_detect_cls_T_1 = cnt_in_detect_cls == 3'h2; // @[control.scala 100:95]
  wire [2:0] _cnt_in_detect_cls_T_3 = cnt_in_detect_cls + 3'h1; // @[control.scala 100:148]
  wire  _layer_finish_T_3 = _conv_cnt_in_c2f_T_3 & conv_finish; // @[control.scala 104:85]
  wire  _layer_finish_T_5 = _cnt_in_sppf_T_1 & conv_finish; // @[control.scala 105:74]
  wire  _layer_finish_T_7 = _cnt_in_detect_box_T_1 & conv_finish; // @[control.scala 106:92]
  wire  _layer_finish_T_9 = _cnt_in_detect_cls_T_1 & conv_finish; // @[control.scala 107:92]
  wire  _layer_finish_T_11 = current_layer_is_detect_box ? _layer_finish_T_7 : current_layer_is_detect_cls &
    _layer_finish_T_9; // @[Mux.scala 101:16]
  wire  _layer_finish_T_12 = current_layer_is_sppf ? _layer_finish_T_5 : _layer_finish_T_11; // @[Mux.scala 101:16]
  wire  _layer_finish_T_13 = current_layer_is_c2f ? _layer_finish_T_3 : _layer_finish_T_12; // @[Mux.scala 101:16]
  wire  layer_finish = current_layer_is_conv ? conv_finish : _layer_finish_T_13; // @[Mux.scala 101:16]
  wire [4:0] _current_layer_T_2 = current_layer + 5'h1; // @[control.scala 109:107]
  reg [15:0] conv_scale; // @[control.scala 112:28]
  reg [3:0] conv_shift; // @[control.scala 113:29]
  reg [7:0] zp_in; // @[control.scala 114:24]
  reg [7:0] zp_out; // @[control.scala 115:25]
  reg [7:0] zp_act; // @[control.scala 116:25]
  reg [31:0] scale_B_act; // @[control.scala 117:30]
  reg [31:0] scale_A_act; // @[control.scala 118:30]
  wire [31:0] reg_scale_shift = {12'h0,conv_shift,conv_scale}; // @[Cat.scala 33:92]
  wire  p_is_1 = current_layer_is_conv | current_layer_is_c2f & (conv_cnt_in_c2f > 5'h0 & conv_cnt_in_c2f <
    _conv_cnt_in_c2f_T_2) | current_layer_is_detect_box & cnt_in_detect_box < 3'h2 | current_layer_is_detect_cls &
    cnt_in_detect_cls < 3'h2; // @[control.scala 269:223]
  wire  k_is_1 = ~p_is_1; // @[control.scala 272:18]
  wire  kernal = ~k_is_1; // @[control.scala 273:15]
  wire [31:0] reg_zp_out_in = {7'h0,kernal,zp_act,zp_out,zp_in}; // @[Cat.scala 33:92]
  wire [31:0] reg_linebuffer_sel = {19'h0,current_layer_sel,10'h0}; // @[Cat.scala 33:92]
  wire [19:0] fm_size_define_0 = 10'h280 * 10'h280; // @[control.scala 128:112]
  wire [17:0] fm_size_define_1 = 9'h140 * 9'h140; // @[control.scala 128:112]
  wire [15:0] fm_size_define_2 = 8'ha0 * 8'ha0; // @[control.scala 128:112]
  wire [13:0] fm_size_define_4 = 7'h50 * 7'h50; // @[control.scala 128:112]
  wire [11:0] fm_size_define_6 = 6'h28 * 6'h28; // @[control.scala 128:112]
  wire [9:0] fm_size_define_8 = 5'h14 * 5'h14; // @[control.scala 128:112]
  wire [4:0] _fm_col_T = cur_layer_sel_21 ? 5'h14 : 5'h0; // @[Mux.scala 101:16]
  wire [5:0] _fm_col_T_1 = cur_layer_sel_20 ? 6'h28 : {{1'd0}, _fm_col_T}; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_2 = cur_layer_sel_19 ? 7'h50 : {{1'd0}, _fm_col_T_1}; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_3 = cur_layer_sel_18 ? 7'h14 : _fm_col_T_2; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_4 = cur_layer_sel_17 ? 7'h28 : _fm_col_T_3; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_5 = cur_layer_sel_16 ? 7'h50 : _fm_col_T_4; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_6 = cur_layer_sel_15 ? 7'h14 : _fm_col_T_5; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_7 = cur_layer_sel_14 ? 7'h28 : _fm_col_T_6; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_8 = cur_layer_sel_13 ? 7'h28 : _fm_col_T_7; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_9 = cur_layer_sel_12 ? 7'h50 : _fm_col_T_8; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_10 = cur_layer_sel_11 ? 7'h50 : _fm_col_T_9; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_11 = cur_layer_sel_10 ? 7'h28 : _fm_col_T_10; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_12 = cur_layer_sel_9 ? 7'h14 : _fm_col_T_11; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_13 = cur_layer_sel_8 ? 7'h14 : _fm_col_T_12; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_14 = cur_layer_sel_7 ? 7'h28 : _fm_col_T_13; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_15 = cur_layer_sel_6 ? 7'h28 : _fm_col_T_14; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_16 = cur_layer_sel_5 ? 7'h50 : _fm_col_T_15; // @[Mux.scala 101:16]
  wire [6:0] _fm_col_T_17 = cur_layer_sel_4 ? 7'h50 : _fm_col_T_16; // @[Mux.scala 101:16]
  wire [7:0] _fm_col_T_18 = cur_layer_sel_3 ? 8'ha0 : {{1'd0}, _fm_col_T_17}; // @[Mux.scala 101:16]
  wire [7:0] _fm_col_T_19 = cur_layer_sel_2 ? 8'ha0 : _fm_col_T_18; // @[Mux.scala 101:16]
  wire [8:0] _fm_col_T_20 = cur_layer_sel_1 ? 9'h140 : {{1'd0}, _fm_col_T_19}; // @[Mux.scala 101:16]
  wire [9:0] fm_col = cur_layer_sel_0 ? 10'h280 : {{1'd0}, _fm_col_T_20}; // @[Mux.scala 101:16]
  wire [9:0] _fm_size_T = cur_layer_sel_21 ? fm_size_define_8 : 10'h0; // @[Mux.scala 101:16]
  wire [11:0] _fm_size_T_1 = cur_layer_sel_20 ? fm_size_define_6 : {{2'd0}, _fm_size_T}; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_2 = cur_layer_sel_19 ? fm_size_define_4 : {{2'd0}, _fm_size_T_1}; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_3 = cur_layer_sel_18 ? {{4'd0}, fm_size_define_8} : _fm_size_T_2; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_4 = cur_layer_sel_17 ? {{2'd0}, fm_size_define_6} : _fm_size_T_3; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_5 = cur_layer_sel_16 ? fm_size_define_4 : _fm_size_T_4; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_6 = cur_layer_sel_15 ? {{4'd0}, fm_size_define_8} : _fm_size_T_5; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_7 = cur_layer_sel_14 ? {{2'd0}, fm_size_define_6} : _fm_size_T_6; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_8 = cur_layer_sel_13 ? {{2'd0}, fm_size_define_6} : _fm_size_T_7; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_9 = cur_layer_sel_12 ? fm_size_define_4 : _fm_size_T_8; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_10 = cur_layer_sel_11 ? fm_size_define_4 : _fm_size_T_9; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_11 = cur_layer_sel_10 ? {{2'd0}, fm_size_define_6} : _fm_size_T_10; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_12 = cur_layer_sel_9 ? {{4'd0}, fm_size_define_8} : _fm_size_T_11; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_13 = cur_layer_sel_8 ? {{4'd0}, fm_size_define_8} : _fm_size_T_12; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_14 = cur_layer_sel_7 ? {{2'd0}, fm_size_define_6} : _fm_size_T_13; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_15 = cur_layer_sel_6 ? {{2'd0}, fm_size_define_6} : _fm_size_T_14; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_16 = cur_layer_sel_5 ? fm_size_define_4 : _fm_size_T_15; // @[Mux.scala 101:16]
  wire [13:0] _fm_size_T_17 = cur_layer_sel_4 ? fm_size_define_4 : _fm_size_T_16; // @[Mux.scala 101:16]
  wire [15:0] _fm_size_T_18 = cur_layer_sel_3 ? fm_size_define_2 : {{2'd0}, _fm_size_T_17}; // @[Mux.scala 101:16]
  wire [15:0] _fm_size_T_19 = cur_layer_sel_2 ? fm_size_define_2 : _fm_size_T_18; // @[Mux.scala 101:16]
  wire [17:0] _fm_size_T_20 = cur_layer_sel_1 ? fm_size_define_1 : {{2'd0}, _fm_size_T_19}; // @[Mux.scala 101:16]
  wire [19:0] _fm_size_T_21 = cur_layer_sel_0 ? fm_size_define_0 : {{2'd0}, _fm_size_T_20}; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_2 = cur_layer_sel_19 ? 6'h2e : _fm_col_T_1; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_3 = cur_layer_sel_18 ? 6'h14 : _fm_div_T_2; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_4 = cur_layer_sel_17 ? 6'h28 : _fm_div_T_3; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_5 = cur_layer_sel_16 ? 6'h2e : _fm_div_T_4; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_6 = cur_layer_sel_15 ? 6'h14 : _fm_div_T_5; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_7 = cur_layer_sel_14 ? 6'h28 : _fm_div_T_6; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_8 = cur_layer_sel_13 ? 6'h28 : _fm_div_T_7; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_9 = cur_layer_sel_12 ? 6'h2e : _fm_div_T_8; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_10 = cur_layer_sel_11 ? 6'h2e : _fm_div_T_9; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_11 = cur_layer_sel_10 ? 6'h28 : _fm_div_T_10; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_12 = cur_layer_sel_9 ? 6'h14 : _fm_div_T_11; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_13 = cur_layer_sel_8 ? 6'h14 : _fm_div_T_12; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_14 = cur_layer_sel_7 ? 6'h28 : _fm_div_T_13; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_15 = cur_layer_sel_6 ? 6'h28 : _fm_div_T_14; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_16 = cur_layer_sel_5 ? 6'h2e : _fm_div_T_15; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_17 = cur_layer_sel_4 ? 6'h2e : _fm_div_T_16; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_18 = cur_layer_sel_3 ? 6'h18 : _fm_div_T_17; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_19 = cur_layer_sel_2 ? 6'h17 : _fm_div_T_18; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_T_20 = cur_layer_sel_1 ? 6'ha : _fm_div_T_19; // @[Mux.scala 101:16]
  wire [5:0] fm_div = cur_layer_sel_0 ? 6'h4 : _fm_div_T_20; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_2 = cur_layer_sel_19 ? 2'h2 : {{1'd0}, _current_layer_repeats_T_1}; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_3 = cur_layer_sel_18 ? 2'h1 : _fm_div_cnt_T_2; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_4 = cur_layer_sel_17 ? 2'h1 : _fm_div_cnt_T_3; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_5 = cur_layer_sel_16 ? 2'h2 : _fm_div_cnt_T_4; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_6 = cur_layer_sel_15 ? 2'h1 : _fm_div_cnt_T_5; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_7 = cur_layer_sel_14 ? 2'h1 : _fm_div_cnt_T_6; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_8 = cur_layer_sel_13 ? 2'h1 : _fm_div_cnt_T_7; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_9 = cur_layer_sel_12 ? 2'h2 : _fm_div_cnt_T_8; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_10 = cur_layer_sel_11 ? 2'h2 : _fm_div_cnt_T_9; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_11 = cur_layer_sel_10 ? 2'h1 : _fm_div_cnt_T_10; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_12 = cur_layer_sel_9 ? 2'h1 : _fm_div_cnt_T_11; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_13 = cur_layer_sel_8 ? 2'h1 : _fm_div_cnt_T_12; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_14 = cur_layer_sel_7 ? 2'h1 : _fm_div_cnt_T_13; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_15 = cur_layer_sel_6 ? 2'h1 : _fm_div_cnt_T_14; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_16 = cur_layer_sel_5 ? 2'h2 : _fm_div_cnt_T_15; // @[Mux.scala 101:16]
  wire [1:0] _fm_div_cnt_T_17 = cur_layer_sel_4 ? 2'h2 : _fm_div_cnt_T_16; // @[Mux.scala 101:16]
  wire [2:0] _fm_div_cnt_T_18 = cur_layer_sel_3 ? 3'h7 : {{1'd0}, _fm_div_cnt_T_17}; // @[Mux.scala 101:16]
  wire [2:0] _fm_div_cnt_T_19 = cur_layer_sel_2 ? 3'h7 : _fm_div_cnt_T_18; // @[Mux.scala 101:16]
  wire [5:0] _fm_div_cnt_T_20 = cur_layer_sel_1 ? 6'h20 : {{3'd0}, _fm_div_cnt_T_19}; // @[Mux.scala 101:16]
  wire [7:0] fm_div_cnt = cur_layer_sel_0 ? 8'ha0 : {{2'd0}, _fm_div_cnt_T_20}; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_2 = cur_layer_sel_19 ? 6'h22 : 6'h0; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_3 = cur_layer_sel_18 ? 6'h0 : _fm_res_T_2; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_4 = cur_layer_sel_17 ? 6'h0 : _fm_res_T_3; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_5 = cur_layer_sel_16 ? 6'h22 : _fm_res_T_4; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_6 = cur_layer_sel_15 ? 6'h0 : _fm_res_T_5; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_7 = cur_layer_sel_14 ? 6'h0 : _fm_res_T_6; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_8 = cur_layer_sel_13 ? 6'h0 : _fm_res_T_7; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_9 = cur_layer_sel_12 ? 6'h22 : _fm_res_T_8; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_10 = cur_layer_sel_11 ? 6'h22 : _fm_res_T_9; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_11 = cur_layer_sel_10 ? 6'h0 : _fm_res_T_10; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_12 = cur_layer_sel_9 ? 6'h0 : _fm_res_T_11; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_13 = cur_layer_sel_8 ? 6'h0 : _fm_res_T_12; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_14 = cur_layer_sel_7 ? 6'h0 : _fm_res_T_13; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_15 = cur_layer_sel_6 ? 6'h0 : _fm_res_T_14; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_16 = cur_layer_sel_5 ? 6'h22 : _fm_res_T_15; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_17 = cur_layer_sel_4 ? 6'h22 : _fm_res_T_16; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_18 = cur_layer_sel_3 ? 6'h10 : _fm_res_T_17; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_19 = cur_layer_sel_2 ? 6'h16 : _fm_res_T_18; // @[Mux.scala 101:16]
  wire [5:0] _fm_res_T_20 = cur_layer_sel_1 ? 6'ha : _fm_res_T_19; // @[Mux.scala 101:16]
  wire [5:0] fm_res = cur_layer_sel_0 ? 6'h4 : _fm_res_T_20; // @[Mux.scala 101:16]
  reg [31:0] reg_t_0; // @[control.scala 160:37]
  reg [31:0] reg_t_1; // @[control.scala 160:37]
  reg [31:0] reg_t_2; // @[control.scala 160:37]
  reg [31:0] reg_t_3; // @[control.scala 160:37]
  reg [31:0] reg_t_4; // @[control.scala 160:37]
  reg [31:0] reg_t_5; // @[control.scala 160:37]
  reg [31:0] reg_t_6; // @[control.scala 160:37]
  reg [31:0] reg_t_7; // @[control.scala 160:37]
  reg [31:0] reg_t_8; // @[control.scala 160:37]
  reg [31:0] reg_t_9; // @[control.scala 160:37]
  reg [31:0] reg_t_10; // @[control.scala 160:37]
  reg [31:0] reg_static; // @[control.scala 161:29]
  reg [31:0] reg_task; // @[control.scala 162:27]
  reg [4:0] cnt_t; // @[control.scala 163:24]
  wire  cnt_t_is_5 = cnt_t == 5'h5; // @[control.scala 165:25]
  reg [31:0] wgt_addr_send; // @[control.scala 178:32]
  reg [15:0] wgt_addr_read; // @[control.scala 179:32]
  reg [15:0] wgt_addr_read_t; // @[control.scala 180:34]
  reg [15:0] bia_addr_read; // @[control.scala 181:32]
  reg  last_buf_sel; // @[control.scala 182:31]
  reg [12:0] iter_ifm_pre; // @[control.scala 192:31]
  reg [12:0] iter_ofm_pre; // @[control.scala 194:31]
  reg [12:0] iter_div_pre; // @[control.scala 195:31]
  reg [12:0] iter_ifm_post; // @[control.scala 196:32]
  reg [12:0] iter_ofm_post; // @[control.scala 197:32]
  reg [12:0] iter_div_post; // @[control.scala 198:32]
  wire  _c2f_cout_T = conv_cnt_in_c2f == 5'h0; // @[control.scala 221:38]
  wire [9:0] current_layer_cout = {{1'd0}, _current_layer_cout_T_21}; // @[control.scala 53:34 64:24]
  wire [9:0] _c2f_cout_T_5 = {{1'd0}, current_layer_cout[9:1]}; // @[control.scala 221:138]
  wire [9:0] _c2f_cout_T_6 = conv_cnt_in_c2f == 5'h0 | _conv_cnt_in_c2f_T_3 ? current_layer_cout : _c2f_cout_T_5; // @[control.scala 221:20]
  wire [15:0] c2f_cout = {{6'd0}, _c2f_cout_T_6}; // @[control.scala 212:24 221:14]
  wire  _sppf_cout_T = cnt_in_sppf == 3'h0; // @[control.scala 223:31]
  wire [9:0] current_layer_cin = {{1'd0}, _current_layer_cin_T_21}; // @[control.scala 54:33 65:23]
  wire [9:0] _sppf_cout_T_2 = cnt_in_sppf == 3'h0 ? {{1'd0}, current_layer_cin[9:1]} : current_layer_cout; // @[control.scala 223:19]
  wire [15:0] sppf_cout = {{6'd0}, _sppf_cout_T_2}; // @[control.scala 214:25 223:14]
  wire  _box_cout_T = ~current_layer_is_detect_box; // @[control.scala 225:47]
  wire [9:0] _box_cout_T_1 = ~current_layer_is_detect_box ? 10'h40 : current_layer_cout; // @[control.scala 225:19]
  wire [15:0] box_cout = {{6'd0}, _box_cout_T_1}; // @[control.scala 216:24 225:14]
  wire  _cls_cout_T = ~current_layer_is_detect_cls; // @[control.scala 227:47]
  wire [9:0] _cls_cout_T_1 = ~current_layer_is_detect_cls ? 10'h50 : current_layer_cout; // @[control.scala 227:19]
  wire [15:0] cls_cout = {{6'd0}, _cls_cout_T_1}; // @[control.scala 218:24 227:14]
  wire [15:0] _cout_T_4 = current_layer_is_detect_cls ? cls_cout : {{6'd0}, current_layer_cout}; // @[Mux.scala 101:16]
  wire [15:0] _cout_T_5 = current_layer_is_detect_box ? box_cout : _cout_T_4; // @[Mux.scala 101:16]
  wire [15:0] _cout_T_6 = current_layer_is_sppf ? sppf_cout : _cout_T_5; // @[Mux.scala 101:16]
  wire [15:0] cout = current_layer_is_c2f ? c2f_cout : _cout_T_6; // @[Mux.scala 101:16]
  wire [12:0] ofm_batch = {{11'd0}, cout[4:3]}; // @[control.scala 188:25 234:14]
  wire [12:0] iter_ofm_post_t = ofm_batch - iter_ofm_post; // @[control.scala 204:34]
  wire [12:0] _GEN_2833 = {{5'd0}, fm_div_cnt}; // @[control.scala 205:35]
  wire [12:0] _iter_div_post_t_T_1 = _GEN_2833 - iter_div_post; // @[control.scala 205:35]
  wire [2:0] _c2f_cin_T_6 = current_layer_repeats + 3'h2; // @[control.scala 220:180]
  wire [9:0] _c2f_cin_T_7 = {{1'd0}, current_layer_cin[9:1]}; // @[control.scala 220:208]
  wire [12:0] _c2f_cin_T_8 = _c2f_cin_T_6 * _c2f_cin_T_7; // @[control.scala 220:187]
  wire [12:0] _c2f_cin_T_9 = _conv_cnt_in_c2f_T_3 ? _c2f_cin_T_8 : {{3'd0}, _c2f_cin_T_7}; // @[Mux.scala 101:16]
  wire [12:0] _c2f_cin_T_10 = _c2f_cout_T ? {{3'd0}, current_layer_cin} : _c2f_cin_T_9; // @[Mux.scala 101:16]
  wire [15:0] c2f_cin = {{3'd0}, _c2f_cin_T_10}; // @[control.scala 213:23 220:13]
  wire [10:0] _sppf_cin_T_1 = {current_layer_cin, 1'h0}; // @[control.scala 222:72]
  wire [10:0] _sppf_cin_T_2 = _sppf_cout_T ? {{1'd0}, current_layer_cin} : _sppf_cin_T_1; // @[control.scala 222:18]
  wire [15:0] sppf_cin = {{5'd0}, _sppf_cin_T_2}; // @[control.scala 215:24 222:13]
  wire [9:0] _box_cin_T_1 = _box_cout_T ? current_layer_cin : 10'h40; // @[control.scala 224:18]
  wire [15:0] box_cin = {{6'd0}, _box_cin_T_1}; // @[control.scala 217:23 224:13]
  wire [9:0] _cls_cin_T_1 = _cls_cout_T ? current_layer_cin : 10'h50; // @[control.scala 226:18]
  wire [15:0] cls_cin = {{6'd0}, _cls_cin_T_1}; // @[control.scala 219:23 226:13]
  wire [15:0] _cin_T_4 = current_layer_is_detect_cls ? cls_cin : {{6'd0}, current_layer_cin}; // @[Mux.scala 101:16]
  wire [15:0] _cin_T_5 = current_layer_is_detect_box ? box_cin : _cin_T_4; // @[Mux.scala 101:16]
  wire [15:0] _cin_T_6 = current_layer_is_sppf ? sppf_cin : _cin_T_5; // @[Mux.scala 101:16]
  wire [15:0] cin = current_layer_is_c2f ? c2f_cin : _cin_T_6; // @[Mux.scala 101:16]
  wire [12:0] ifm_batch = {{11'd0}, cin[4:3]}; // @[control.scala 189:25 235:14]
  wire [12:0] _iter_ifm_post_t_T_1 = ifm_batch - iter_ifm_post; // @[control.scala 206:34]
  wire [12:0] _iter_div_pre_t_T_1 = _GEN_2833 - iter_div_pre; // @[control.scala 207:34]
  wire [12:0] iter_ifm_pre_t = ifm_batch - iter_ifm_pre; // @[control.scala 208:33]
  wire  _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_1 = current_layer_is_detect_box & cnt_in_detect_box != 3'h0; // @[control.scala 260:142]
  wire  _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_3 = current_layer_is_detect_cls & cnt_in_detect_cls != 3'h0; // @[control.scala 260:238]
  wire  ifm_batch_is_exactly_divided_by_WEIGHT_LEN_temp = cur_layer_sel_0 | (cur_layer_sel_1 | (cur_layer_sel_2 | (
    cur_layer_sel_3 | (cur_layer_sel_4 | (cur_layer_sel_5 | (cur_layer_sel_6 | (cur_layer_sel_7 | (cur_layer_sel_8 | (
    cur_layer_sel_9 | (cur_layer_sel_10 | (cur_layer_sel_11 | (cur_layer_sel_12 | (cur_layer_sel_13 | (cur_layer_sel_14
     | (cur_layer_sel_15 | (cur_layer_sel_16 | (cur_layer_sel_17 | (cur_layer_sel_18 | (cur_layer_sel_19 | (
    cur_layer_sel_20 | cur_layer_sel_21)))))))))))))))))))); // @[Mux.scala 101:16]
  wire  _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_4 = _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_3 ? 1'h0 :
    ifm_batch_is_exactly_divided_by_WEIGHT_LEN_temp; // @[Mux.scala 101:16]
  wire  ifm_batch_is_exactly_divided_by_WEIGHT_LEN = _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_1 |
    _ifm_batch_is_exactly_divided_by_WEIGHT_LEN_T_4; // @[Mux.scala 101:16]
  wire  _skip_act_T_1 = current_layer_is_detect_box & _cnt_in_detect_box_T_1; // @[control.scala 265:46]
  wire  _skip_act_T_3 = current_layer_is_detect_cls & _cnt_in_detect_cls_T_1; // @[control.scala 265:135]
  wire  skip_act = current_layer_is_detect_box & _cnt_in_detect_box_T_1 | current_layer_is_detect_cls &
    _cnt_in_detect_cls_T_1; // @[control.scala 265:103]
  reg [2:0] weight_sel; // @[control.scala 274:27]
  wire [25:0] _weight_len_limit_T = ifm_batch * ofm_batch; // @[control.scala 276:43]
  wire [25:0] weight_len_limit = _weight_len_limit_T <= 26'h80 ? _weight_len_limit_T : 26'h80; // @[control.scala 276:31]
  wire [25:0] _weight_len_T = ifm_batch_is_exactly_divided_by_WEIGHT_LEN ? weight_len_limit : {{13'd0}, ifm_batch}; // @[control.scala 277:20]
  wire [5:0] _upsample_start_batch_T = cur_layer_sel_21 ? 6'h20 : 6'h0; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_1 = cur_layer_sel_20 ? 6'h10 : _upsample_start_batch_T; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_2 = cur_layer_sel_19 ? 6'h8 : _upsample_start_batch_T_1; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_3 = cur_layer_sel_18 ? 6'h20 : _upsample_start_batch_T_2; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_4 = cur_layer_sel_17 ? 6'h10 : _upsample_start_batch_T_3; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_5 = cur_layer_sel_16 ? 6'h8 : _upsample_start_batch_T_4; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_6 = cur_layer_sel_15 ? 6'h30 : _upsample_start_batch_T_5; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_7 = cur_layer_sel_14 ? 6'h10 : _upsample_start_batch_T_6; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_8 = cur_layer_sel_13 ? 6'h18 : _upsample_start_batch_T_7; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_9 = cur_layer_sel_12 ? 6'h8 : _upsample_start_batch_T_8; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_10 = cur_layer_sel_11 ? 6'h8 : _upsample_start_batch_T_9; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_11 = cur_layer_sel_10 ? 6'h10 : _upsample_start_batch_T_10; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_12 = cur_layer_sel_9 ? 6'h20 : _upsample_start_batch_T_11; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_13 = cur_layer_sel_8 ? 6'h20 : _upsample_start_batch_T_12; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_14 = cur_layer_sel_7 ? 6'h10 : _upsample_start_batch_T_13; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_15 = cur_layer_sel_6 ? 6'h10 : _upsample_start_batch_T_14; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_16 = cur_layer_sel_5 ? 6'h8 : _upsample_start_batch_T_15; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_17 = cur_layer_sel_4 ? 6'h8 : _upsample_start_batch_T_16; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_18 = cur_layer_sel_3 ? 6'h4 : _upsample_start_batch_T_17; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_19 = cur_layer_sel_2 ? 6'h4 : _upsample_start_batch_T_18; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_20 = cur_layer_sel_1 ? 6'h2 : _upsample_start_batch_T_19; // @[Mux.scala 101:16]
  wire [5:0] _upsample_start_batch_T_21 = cur_layer_sel_0 ? 6'h1 : _upsample_start_batch_T_20; // @[Mux.scala 101:16]
  wire  _upsample_en_T_1 = current_layer_is_c2f & _c2f_cout_T; // @[control.scala 283:39]
  wire [9:0] upsample_start_batch = {{4'd0}, _upsample_start_batch_T_21}; // @[control.scala 279:36 281:26]
  wire [12:0] _GEN_2839 = {{3'd0}, upsample_start_batch}; // @[control.scala 283:82]
  wire  upsample_en = current_layer_is_c2f & _c2f_cout_T & iter_ifm_pre >= _GEN_2839; // @[control.scala 283:66]
  wire [13:0] _c2f_size_half_T = cur_layer_sel_21 ? 14'h3e80 : 14'h0; // @[Mux.scala 101:16]
  wire [15:0] _c2f_size_half_T_1 = cur_layer_sel_20 ? 16'hfa00 : {{2'd0}, _c2f_size_half_T}; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_2 = cur_layer_sel_19 ? 18'h3e800 : {{2'd0}, _c2f_size_half_T_1}; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_3 = cur_layer_sel_18 ? 18'h3200 : _c2f_size_half_T_2; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_4 = cur_layer_sel_17 ? 18'hc800 : _c2f_size_half_T_3; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_5 = cur_layer_sel_16 ? 18'h32000 : _c2f_size_half_T_4; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_6 = cur_layer_sel_15 ? 18'hc800 : _c2f_size_half_T_5; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_7 = cur_layer_sel_14 ? 18'h19000 : _c2f_size_half_T_6; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_8 = cur_layer_sel_13 ? 18'h19000 : _c2f_size_half_T_7; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_9 = cur_layer_sel_12 ? 18'h32000 : _c2f_size_half_T_8; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_10 = cur_layer_sel_11 ? 18'h32000 : _c2f_size_half_T_9; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_11 = cur_layer_sel_10 ? 18'h19000 : _c2f_size_half_T_10; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_12 = cur_layer_sel_9 ? 18'hc800 : _c2f_size_half_T_11; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_13 = cur_layer_sel_8 ? 18'hc800 : _c2f_size_half_T_12; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_14 = cur_layer_sel_7 ? 18'h32000 : _c2f_size_half_T_13; // @[Mux.scala 101:16]
  wire [17:0] _c2f_size_half_T_15 = cur_layer_sel_6 ? 18'h19000 : _c2f_size_half_T_14; // @[Mux.scala 101:16]
  wire [18:0] _c2f_size_half_T_16 = cur_layer_sel_5 ? 19'h64000 : {{1'd0}, _c2f_size_half_T_15}; // @[Mux.scala 101:16]
  wire [18:0] _c2f_size_half_T_17 = cur_layer_sel_4 ? 19'h32000 : _c2f_size_half_T_16; // @[Mux.scala 101:16]
  wire [19:0] _c2f_size_half_T_18 = cur_layer_sel_3 ? 20'hc8000 : {{1'd0}, _c2f_size_half_T_17}; // @[Mux.scala 101:16]
  wire [19:0] _c2f_size_half_T_19 = cur_layer_sel_2 ? 20'h64000 : _c2f_size_half_T_18; // @[Mux.scala 101:16]
  wire [20:0] _c2f_size_half_T_20 = cur_layer_sel_1 ? 21'h190000 : {{1'd0}, _c2f_size_half_T_19}; // @[Mux.scala 101:16]
  wire [21:0] _c2f_size_half_T_21 = cur_layer_sel_0 ? 22'h320000 : {{1'd0}, _c2f_size_half_T_20}; // @[Mux.scala 101:16]
  wire  pool_en = current_layer_is_sppf & _sppf_cout_T; // @[control.scala 289:38]
  reg [1:0] pool_cnt; // @[control.scala 290:27]
  wire  _pool_addr_base_T = pool_cnt == 2'h0; // @[control.scala 292:52]
  wire  _pool_addr_base_T_1 = pool_cnt == 2'h1; // @[control.scala 292:90]
  wire  _pool_addr_base_T_2 = pool_cnt == 2'h2; // @[control.scala 292:128]
  wire  _pool_addr_base_T_3 = pool_cnt == 2'h3; // @[control.scala 292:166]
  wire [29:0] _pool_addr_base_T_4 = _pool_addr_base_T_3 ? 30'h20ca5800 : 30'h0; // @[Mux.scala 101:16]
  wire [29:0] _pool_addr_base_T_5 = _pool_addr_base_T_2 ? 30'h20c99000 : _pool_addr_base_T_4; // @[Mux.scala 101:16]
  wire [29:0] _pool_addr_base_T_6 = _pool_addr_base_T_1 ? 30'h20c8c800 : _pool_addr_base_T_5; // @[Mux.scala 101:16]
  wire [29:0] _pool_addr_base_T_7 = _pool_addr_base_T ? 30'h20c80000 : _pool_addr_base_T_6; // @[Mux.scala 101:16]
  reg  bottleneck_transfer; // @[control.scala 295:38]
  reg  bottleneck_ready; // @[control.scala 296:35]
  wire  _bottleneck_en_T_1 = conv_cnt_in_c2f != 5'h0; // @[control.scala 297:79]
  wire  _bottleneck_en_T_5 = conv_cnt_in_c2f != _conv_cnt_in_c2f_T_2; // @[control.scala 297:108]
  wire  _bottleneck_en_T_8 = ~conv_cnt_in_c2f[0]; // @[control.scala 297:163]
  wire  bottleneck_en = c2f_shortcut & current_layer_is_c2f & conv_cnt_in_c2f != 5'h0 & conv_cnt_in_c2f !=
    _conv_cnt_in_c2f_T_2 & ~conv_cnt_in_c2f[0]; // @[control.scala 297:140]
  reg [1:0] cnt_detect_cls; // @[control.scala 299:33]
  reg  current_layer_is_detect_cls_next; // @[control.scala 300:51]
  wire [1:0] _cnt_detect_cls_T_4 = cnt_detect_cls + 2'h1; // @[control.scala 301:172]
  wire  _ofm_write_disable_T = _iter_ifm_post_t_T_1 == 13'h1; // @[control.scala 304:44]
  wire  _ofm_write_disable_T_1 = ~bottleneck_ready; // @[control.scala 304:56]
  wire  ofm_write_disable = ~(_iter_ifm_post_t_T_1 == 13'h1 & ~bottleneck_ready); // @[control.scala 304:26]
  wire [31:0] _reg_t_8_T_1 = {8'h0,ifm_batch[3:0],cnt_detect_cls,ofm_write_disable,_skip_act_T_3,4'h0,pool_cnt,fm_col}; // @[Cat.scala 33:92]
  reg [31:0] iter_div_prexfm_div_col; // @[control.scala 316:41]
  reg [31:0] fm_row_fm_res_t1xfm_col; // @[control.scala 319:41]
  reg [31:0] fm_row_fm_resxfm_col; // @[control.scala 320:38]
  wire [15:0] _fm_div_col_T = fm_div * fm_col; // @[control.scala 324:26]
  wire [5:0] fm_div_t2 = fm_div + 6'h2; // @[control.scala 325:25]
  wire [5:0] fm_div_t1 = fm_div + 6'h1; // @[control.scala 326:25]
  wire [5:0] fm_res_t1 = fm_res + 6'h1; // @[control.scala 328:25]
  wire [14:0] fm_div_col = _fm_div_col_T[14:0]; // @[control.scala 314:24 324:16]
  wire [27:0] _iter_div_prexfm_div_col_T = iter_div_pre * fm_div_col; // @[control.scala 332:44]
  wire [9:0] _GEN_2841 = {{4'd0}, fm_res_t1}; // @[control.scala 334:38]
  wire [9:0] _fm_row_fm_res_t1xfm_col_T_1 = fm_col - _GEN_2841; // @[control.scala 334:38]
  wire [19:0] _fm_row_fm_res_t1xfm_col_T_2 = _fm_row_fm_res_t1xfm_col_T_1 * fm_col; // @[control.scala 334:50]
  wire [9:0] _GEN_2842 = {{4'd0}, fm_res}; // @[control.scala 335:35]
  wire [9:0] _fm_row_fm_resxfm_col_T_1 = fm_col - _GEN_2842; // @[control.scala 335:35]
  wire [19:0] _fm_row_fm_resxfm_col_T_2 = _fm_row_fm_resxfm_col_T_1 * fm_col; // @[control.scala 335:44]
  wire [18:0] fm_size = _fm_size_T_21[18:0]; // @[control.scala 131:23 136:13]
  wire [18:0] fm_size_output = current_layer_is_conv ? {{2'd0}, fm_size[18:2]} : fm_size; // @[control.scala 347:26]
  wire [9:0] fm_col_output = current_layer_is_conv ? {{1'd0}, fm_col[9:1]} : fm_col; // @[control.scala 348:25]
  wire  _fm_div_output_T = current_layer_is_conv & p_is_1; // @[control.scala 349:32]
  wire [5:0] fm_div_output = current_layer_is_conv & p_is_1 ? {{1'd0}, fm_div[5:1]} : fm_div; // @[control.scala 349:25]
  wire [5:0] fm_res_output = _fm_div_output_T ? {{1'd0}, fm_res[5:1]} : fm_res; // @[control.scala 350:25]
  reg [31:0] iter_div_postxfm_col_output; // @[control.scala 352:44]
  reg [31:0] fm_row_res_outputxfm_col_output; // @[control.scala 353:48]
  wire [18:0] _iter_div_postxfm_col_output_T = iter_div_post * fm_div_output; // @[control.scala 354:47]
  wire [28:0] _iter_div_postxfm_col_output_T_1 = _iter_div_postxfm_col_output_T * fm_col_output; // @[control.scala 354:61]
  wire [9:0] _GEN_2843 = {{4'd0}, fm_res_output}; // @[control.scala 355:54]
  wire [9:0] _fm_row_res_outputxfm_col_output_T_1 = fm_col_output - _GEN_2843; // @[control.scala 355:54]
  wire [19:0] _fm_row_res_outputxfm_col_output_T_2 = _fm_row_res_outputxfm_col_output_T_1 * fm_col_output; // @[control.scala 355:69]
  reg  ifm_send_task_enable; // @[control.scala 357:39]
  reg  ofm_recv_task_enable; // @[control.scala 358:39]
  reg  wgt_send_task_enable; // @[control.scala 359:39]
  reg [31:0] ifm_addr_fmbase; // @[control.scala 362:34]
  reg [31:0] ifm_addr_offset; // @[control.scala 363:34]
  reg [31:0] ifm_send_len; // @[control.scala 364:31]
  reg [31:0] ofm_addr_fmbase; // @[control.scala 365:34]
  reg [31:0] ofm_addr_offset; // @[control.scala 366:34]
  reg [31:0] ofm_recv_len; // @[control.scala 367:31]
  reg [31:0] wgt_ddr_base_addr; // @[control.scala 369:36]
  reg [31:0] bia_ddr_base_addr; // @[control.scala 370:36]
  reg  ifm_sel; // @[control.scala 379:24]
  reg [31:0] ifm_addr_t; // @[control.scala 380:29]
  reg [31:0] ifm_addr_send; // @[control.scala 381:32]
  wire [29:0] _ifm_addr_base_T = ifm_sel ? 30'h20320000 : 30'h20000000; // @[control.scala 382:23]
  wire [31:0] ifm_addr_base = {{2'd0}, _ifm_addr_base_T}; // @[control.scala 374:29 382:18]
  wire [31:0] _ifm_ddr_base_addr_t_T_1 = 5'h0 == current_layer ? ifm_addr_base : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_3 = 5'h1 == current_layer ? 32'h207d0000 : _ifm_ddr_base_addr_t_T_1; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_5 = 5'h2 == current_layer ? 32'h20640000 : _ifm_ddr_base_addr_t_T_3; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_7 = 5'h3 == current_layer ? 32'h207d0000 : _ifm_ddr_base_addr_t_T_5; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_9 = 5'h4 == current_layer ? 32'h20640000 : _ifm_ddr_base_addr_t_T_7; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_11 = 5'h5 == current_layer ? 32'h20cb2000 : _ifm_ddr_base_addr_t_T_9; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_13 = 5'h6 == current_layer ? 32'h207d0000 : _ifm_ddr_base_addr_t_T_11; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_15 = 5'h7 == current_layer ? 32'h20d61000 : _ifm_ddr_base_addr_t_T_13; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_17 = 5'h8 == current_layer ? 32'h20640000 : _ifm_ddr_base_addr_t_T_15; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_19 = 5'h9 == current_layer ? 32'h207d0000 : _ifm_ddr_base_addr_t_T_17; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_21 = 5'ha == current_layer ? 32'h20d61000 : _ifm_ddr_base_addr_t_T_19; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_23 = 5'hb == current_layer ? 32'h20cb2000 : _ifm_ddr_base_addr_t_T_21; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_25 = 5'hc == current_layer ? 32'h20db8800 : _ifm_ddr_base_addr_t_T_23; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_27 = 5'hd == current_layer ? 32'h20d16000 : _ifm_ddr_base_addr_t_T_25; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_29 = 5'he == current_layer ? 32'h20e1c800 : _ifm_ddr_base_addr_t_T_27; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_31 = 5'hf == current_layer ? 32'h20d93000 : _ifm_ddr_base_addr_t_T_29; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_33 = 5'h10 == current_layer ? 32'h20db8800 : _ifm_ddr_base_addr_t_T_31; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_35 = 5'h11 == current_layer ? 32'h20e1c800 : _ifm_ddr_base_addr_t_T_33; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_37 = 5'h12 == current_layer ? 32'h20e4e800 : _ifm_ddr_base_addr_t_T_35; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_39 = 5'h13 == current_layer ? 32'h20db8800 : _ifm_ddr_base_addr_t_T_37; // @[Mux.scala 81:58]
  wire [31:0] _ifm_ddr_base_addr_t_T_41 = 5'h14 == current_layer ? 32'h20e1c800 : _ifm_ddr_base_addr_t_T_39; // @[Mux.scala 81:58]
  wire [31:0] ifm_ddr_base_addr_t = 5'h15 == current_layer ? 32'h20e4e800 : _ifm_ddr_base_addr_t_T_41; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_1 = 5'h0 == current_layer ? 30'h207d0000 : 30'h0; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_3 = 5'h1 == current_layer ? 30'h20640000 : _ofm_ddr_base_addr_t_T_1; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_5 = 5'h2 == current_layer ? 30'h207d0000 : _ofm_ddr_base_addr_t_T_3; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_7 = 5'h3 == current_layer ? 30'h20640000 : _ofm_ddr_base_addr_t_T_5; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_9 = 5'h4 == current_layer ? 30'h20cb2000 : _ofm_ddr_base_addr_t_T_7; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_11 = 5'h5 == current_layer ? 30'h207d0000 : _ofm_ddr_base_addr_t_T_9; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_13 = 5'h6 == current_layer ? 30'h20d61000 : _ofm_ddr_base_addr_t_T_11; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_15 = 5'h7 == current_layer ? 30'h20640000 : _ofm_ddr_base_addr_t_T_13; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_17 = 5'h8 == current_layer ? 30'h207d0000 : _ofm_ddr_base_addr_t_T_15; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_19 = 5'h9 == current_layer ? 30'h20d93000 : _ofm_ddr_base_addr_t_T_17; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_21 = 5'ha == current_layer ? 30'h20d16000 : _ofm_ddr_base_addr_t_T_19; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_23 = 5'hb == current_layer ? 30'h20db8800 : _ofm_ddr_base_addr_t_T_21; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_25 = 5'hc == current_layer ? 30'h20d48000 : _ofm_ddr_base_addr_t_T_23; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_27 = 5'hd == current_layer ? 30'h20e1c800 : _ofm_ddr_base_addr_t_T_25; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_29 = 5'he == current_layer ? 30'h20dac000 : _ofm_ddr_base_addr_t_T_27; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_31 = 5'hf == current_layer ? 30'h20e4e800 : _ofm_ddr_base_addr_t_T_29; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_33 = 5'h10 == current_layer ? 30'h20e67800 : _ofm_ddr_base_addr_t_T_31; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_35 = 5'h11 == current_layer ? 30'h20ecb800 : _ofm_ddr_base_addr_t_T_33; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_37 = 5'h12 == current_layer ? 30'h20ee4800 : _ofm_ddr_base_addr_t_T_35; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_39 = 5'h13 == current_layer ? 30'h20eeac00 : _ofm_ddr_base_addr_t_T_37; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_41 = 5'h14 == current_layer ? 30'h20f67c00 : _ofm_ddr_base_addr_t_T_39; // @[Mux.scala 81:58]
  wire [29:0] _ofm_ddr_base_addr_t_T_43 = 5'h15 == current_layer ? 30'h20f87000 : _ofm_ddr_base_addr_t_T_41; // @[Mux.scala 81:58]
  wire [4:0] _cnt_n_in_c2f_T_1 = conv_cnt_in_c2f - 5'h1; // @[control.scala 397:35]
  wire [2:0] cnt_n_in_c2f = _cnt_n_in_c2f_T_1[3:1]; // @[control.scala 396:26 397:17]
  wire [2:0] _ifm_ddr_base_addr_temp_c2f_one_T_4 = cnt_n_in_c2f + 3'h1; // @[control.scala 398:134]
  wire [31:0] c2f_size_half = {{10'd0}, _c2f_size_half_T_21}; // @[control.scala 284:29 286:19]
  wire [34:0] _ifm_ddr_base_addr_temp_c2f_one_T_5 = _ifm_ddr_base_addr_temp_c2f_one_T_4 * c2f_size_half; // @[control.scala 398:141]
  wire [34:0] _ifm_ddr_base_addr_temp_c2f_one_T_7 = 35'h20960000 + _ifm_ddr_base_addr_temp_c2f_one_T_5; // @[control.scala 398:118]
  wire [34:0] _ifm_ddr_base_addr_temp_c2f_one_T_8 = _conv_cnt_in_c2f_T_3 ? 35'h20960000 :
    _ifm_ddr_base_addr_temp_c2f_one_T_7; // @[control.scala 398:42]
  wire [2:0] _ofm_ddr_base_addr_temp_c2f_two_T_2 = cnt_n_in_c2f + 3'h2; // @[control.scala 400:102]
  wire [34:0] _ofm_ddr_base_addr_temp_c2f_two_T_3 = _ofm_ddr_base_addr_temp_c2f_two_T_2 * c2f_size_half; // @[control.scala 400:109]
  wire [34:0] _ofm_ddr_base_addr_temp_c2f_two_T_4 = _c2f_cout_T ? 35'h0 : _ofm_ddr_base_addr_temp_c2f_two_T_3; // @[control.scala 400:57]
  wire [34:0] _ofm_ddr_base_addr_temp_c2f_two_T_6 = 35'h20960000 + _ofm_ddr_base_addr_temp_c2f_two_T_4; // @[control.scala 400:52]
  wire  _ifm_ddr_base_addr_temp_c2f_T_4 = _bottleneck_en_T_1 & _bottleneck_en_T_5; // @[control.scala 401:65]
  wire [31:0] ifm_ddr_base_addr_temp_c2f_one = _ifm_ddr_base_addr_temp_c2f_one_T_8[31:0]; // @[control.scala 394:46 398:36]
  wire [31:0] ifm_ddr_base_addr_temp_c2f = _bottleneck_en_T_1 & _bottleneck_en_T_5 & _bottleneck_en_T_8 ? 32'h20af0000
     : ifm_ddr_base_addr_temp_c2f_one; // @[control.scala 401:38]
  wire [31:0] ofm_ddr_base_addr_temp_c2f_two = _ofm_ddr_base_addr_temp_c2f_two_T_6[31:0]; // @[control.scala 395:46 400:36]
  wire [31:0] ofm_ddr_base_addr_temp_c2f = _ifm_ddr_base_addr_temp_c2f_T_4 & conv_cnt_in_c2f[0] ? 32'h20af0000 :
    ofm_ddr_base_addr_temp_c2f_two; // @[control.scala 402:38]
  wire [29:0] _ifm_ddr_base_addr_temp_sppf_T_3 = _sppf_cout_T ? 30'h207d0000 : 30'h20c80000; // @[Mux.scala 101:16]
  wire [29:0] _ofm_ddr_base_addr_temp_sppf_T_2 = _cnt_in_sppf_T_1 ? 30'h20d93000 : 30'h20c80000; // @[Mux.scala 101:16]
  wire [31:0] pool_addr_base = {{2'd0}, _pool_addr_base_T_7}; // @[control.scala 291:30 292:20]
  wire [31:0] ofm_ddr_base_addr_temp_sppf = _sppf_cout_T ? pool_addr_base : {{2'd0}, _ofm_ddr_base_addr_temp_sppf_T_2}; // @[Mux.scala 101:16]
  wire [31:0] ifm_ddr_base_addr_temp_sppf = {{2'd0}, _ifm_ddr_base_addr_temp_sppf_T_3}; // @[control.scala 392:43 403:33]
  wire [31:0] _ifm_ddr_base_addr_temp_T = current_layer_is_sppf ? ifm_ddr_base_addr_temp_sppf : 32'h20af0000; // @[control.scala 405:88]
  wire [31:0] ifm_ddr_base_addr_temp = current_layer_is_c2f ? ifm_ddr_base_addr_temp_c2f : _ifm_ddr_base_addr_temp_T; // @[control.scala 405:34]
  wire [31:0] _ofm_ddr_base_addr_temp_T = current_layer_is_sppf ? ofm_ddr_base_addr_temp_sppf : 32'h20af0000; // @[control.scala 406:88]
  wire [31:0] ofm_ddr_base_addr_temp = current_layer_is_c2f ? ofm_ddr_base_addr_temp_c2f : _ofm_ddr_base_addr_temp_T; // @[control.scala 406:34]
  wire [31:0] ifm_ddr_base_addr = current_layer_is_conv | _upsample_en_T_1 | pool_en | current_layer_is_detect_cls &
    cnt_in_detect_cls == 3'h0 | current_layer_is_detect_box & cnt_in_detect_box == 3'h0 ? ifm_ddr_base_addr_t :
    ifm_ddr_base_addr_temp; // @[control.scala 408:29]
  wire [31:0] ofm_ddr_base_addr_t = {{2'd0}, _ofm_ddr_base_addr_t_T_43}; // @[control.scala 376:35 385:24]
  wire [31:0] ofm_ddr_base_addr = current_layer_is_conv | current_layer_is_c2f & _conv_cnt_in_c2f_T_3 |
    current_layer_is_sppf & _cnt_in_sppf_T_1 | _skip_act_T_3 | _skip_act_T_1 ? ofm_ddr_base_addr_t :
    ofm_ddr_base_addr_temp; // @[control.scala 409:29]
  reg [31:0] ifm_ddr_base_addr_regnext1; // @[Reg.scala 35:20]
  reg [31:0] ifm_ddr_base_addr_regnext2; // @[Reg.scala 35:20]
  wire [31:0] _ifm_addr_t_T_1 = ifm_addr_fmbase + ifm_addr_offset; // @[control.scala 413:36]
  wire [34:0] _ifm_addr_t_T_2 = {_ifm_addr_t_T_1, 3'h0}; // @[control.scala 413:55]
  wire [31:0] _ifm_addr_send_T = bottleneck_transfer ? ifm_ddr_base_addr_regnext2 : ifm_ddr_base_addr; // @[control.scala 414:25]
  wire [31:0] _ifm_addr_send_T_2 = _ifm_addr_send_T + ifm_addr_t; // @[control.scala 414:92]
  reg [31:0] ofm_addr_t; // @[control.scala 415:29]
  reg [31:0] ofm_addr_recv; // @[control.scala 416:32]
  wire [31:0] _ofm_addr_t_T_1 = ofm_addr_fmbase + ofm_addr_offset; // @[control.scala 417:36]
  wire [34:0] _ofm_addr_t_T_2 = {_ofm_addr_t_T_1, 3'h0}; // @[control.scala 417:55]
  wire [31:0] _ofm_addr_recv_T_1 = ofm_ddr_base_addr + ofm_addr_t; // @[control.scala 418:40]
  reg  resize_load_t; // @[control.scala 420:32]
  reg  first_ofm_recv_stop; // @[control.scala 422:38]
  reg  wgt_ddr_read_en; // @[control.scala 424:32]
  reg [7:0] the_number_of_row_transferred; // @[control.scala 425:46]
  reg [5:0] state; // @[control.scala 436:24]
  wire [4:0] _cnt_t_T_1 = cnt_t + 5'h1; // @[control.scala 449:32]
  wire [4:0] _GEN_2 = cnt_t_is_5 ? 5'h0 : _cnt_t_T_1; // @[control.scala 445:30 446:23 449:23]
  wire [18:0] _reg_t_5_T = {ofm_batch, 6'h0}; // @[control.scala 474:35]
  wire [5:0] _GEN_6 = cnt_t_is_5 ? 6'h3 : state; // @[control.scala 480:30 482:23 436:24]
  wire [31:0] _GEN_7 = cnt_t_is_5 ? 32'h8 : reg_t_0; // @[control.scala 480:30 483:26 160:37]
  wire [2:0] _GEN_8 = ap_done_up ? 3'h4 : 3'h3; // @[control.scala 490:30 491:23 493:23]
  wire [4:0] _reg_t_5_T_1 = 1'h1 * 4'h8; // @[control.scala 499:41]
  wire [8:0] _reg_t_5_T_2 = _reg_t_5_T_1 * 4'h8; // @[control.scala 499:47]
  wire [7:0] _reg_t_5_T_3 = 4'h9 * 4'h8; // @[control.scala 499:61]
  wire [11:0] _reg_t_5_T_4 = _reg_t_5_T_3 * 4'h8; // @[control.scala 499:67]
  wire [7:0] weight_len = _weight_len_T[7:0]; // @[control.scala 275:24 277:15]
  wire [19:0] _reg_t_5_T_5 = _reg_t_5_T_4 * weight_len; // @[control.scala 499:73]
  wire [19:0] _reg_t_5_T_6 = k_is_1 ? {{11'd0}, _reg_t_5_T_2} : _reg_t_5_T_5; // @[control.scala 499:28]
  wire [5:0] _GEN_10 = cnt_t_is_5 ? 6'h6 : state; // @[control.scala 505:30 507:23 436:24]
  wire [31:0] _GEN_11 = cnt_t_is_5 ? 32'h4 : reg_t_0; // @[control.scala 505:30 508:26 160:37]
  wire [31:0] _GEN_12 = cnt_t_is_5 ? reg_scale_shift : reg_t_1; // @[control.scala 505:30 510:26 160:37]
  wire [31:0] _GEN_13 = cnt_t_is_5 ? reg_zp_out_in : reg_t_2; // @[control.scala 505:30 511:26 160:37]
  wire [31:0] _GEN_14 = cnt_t_is_5 ? scale_B_act : reg_t_9; // @[control.scala 505:30 512:26 160:37]
  wire [31:0] _GEN_15 = cnt_t_is_5 ? scale_A_act : reg_t_10; // @[control.scala 505:30 513:27 160:37]
  wire [2:0] _GEN_16 = ap_done_up ? 3'h7 : 3'h6; // @[control.scala 520:30 521:23 523:23]
  wire  _T_9 = iter_ofm_post_t != 13'h1; // @[control.scala 530:34]
  wire  _T_13 = iter_ofm_post_t != 13'h1 | _iter_div_post_t_T_1 != 13'h1 | _iter_ifm_post_t_T_1 != 13'h1; // @[control.scala 530:69]
  wire [3:0] _GEN_18 = iter_ofm_post_t != 13'h1 | _iter_div_post_t_T_1 != 13'h1 | _iter_ifm_post_t_T_1 != 13'h1 ? 4'h8
     : 4'h9; // @[control.scala 530:97 532:23 535:23]
  wire [31:0] _ifm_addr_fmbase_T = iter_ifm_pre * fm_size; // @[control.scala 540:45]
  wire  _T_15 = fm_div_cnt == 8'h1; // @[control.scala 543:29]
  wire [21:0] _ifm_send_len_T = {fm_size, 3'h0}; // @[control.scala 548:41]
  wire  _T_16 = _iter_div_pre_t_T_1 == 13'h1; // @[control.scala 555:45]
  wire [15:0] _ifm_send_len_T_1 = fm_res_t1 * fm_col; // @[control.scala 557:56]
  wire [18:0] _ifm_send_len_T_2 = {_ifm_send_len_T_1, 3'h0}; // @[control.scala 557:66]
  wire  _T_17 = iter_div_pre == 13'h0; // @[control.scala 559:49]
  wire [18:0] _ifm_send_len_T_4 = {_fm_div_col_T, 3'h0}; // @[control.scala 561:63]
  wire [31:0] _GEN_2844 = {{22'd0}, fm_col}; // @[control.scala 564:72]
  wire [31:0] _ifm_addr_offset_T_1 = iter_div_prexfm_div_col - _GEN_2844; // @[control.scala 564:72]
  wire [15:0] _ifm_send_len_T_5 = fm_div_t1 * fm_col; // @[control.scala 565:56]
  wire [18:0] _ifm_send_len_T_6 = {_ifm_send_len_T_5, 3'h0}; // @[control.scala 565:66]
  wire [31:0] _GEN_19 = iter_div_pre == 13'h0 ? 32'h0 : _ifm_addr_offset_T_1; // @[control.scala 559:58 560:45 564:45]
  wire [18:0] _GEN_20 = iter_div_pre == 13'h0 ? _ifm_send_len_T_4 : _ifm_send_len_T_6; // @[control.scala 559:58 561:42 565:42]
  wire [5:0] _GEN_21 = iter_div_pre == 13'h0 ? fm_div : fm_div_t1; // @[control.scala 559:58 562:59 566:59]
  wire [31:0] _GEN_22 = _iter_div_pre_t_T_1 == 13'h1 ? fm_row_fm_res_t1xfm_col : _GEN_19; // @[control.scala 555:54 556:45]
  wire [18:0] _GEN_23 = _iter_div_pre_t_T_1 == 13'h1 ? _ifm_send_len_T_2 : _GEN_20; // @[control.scala 555:54 557:42]
  wire [5:0] _GEN_24 = _iter_div_pre_t_T_1 == 13'h1 ? fm_res_t1 : _GEN_21; // @[control.scala 555:54 558:59]
  wire [31:0] _reg_static_T = reg_linebuffer_sel | 32'h40000; // @[control.scala 568:58]
  wire [31:0] _GEN_25 = p_is_1 ? _GEN_22 : ifm_addr_offset; // @[control.scala 363:34 554:35]
  wire [31:0] _GEN_26 = p_is_1 ? {{13'd0}, _GEN_23} : ifm_send_len; // @[control.scala 364:31 554:35]
  wire [7:0] _GEN_27 = p_is_1 ? {{2'd0}, _GEN_24} : the_number_of_row_transferred; // @[control.scala 554:35 425:46]
  wire [31:0] _GEN_28 = p_is_1 ? _reg_static_T : reg_static; // @[control.scala 161:29 554:35 568:36]
  wire [15:0] _ifm_send_len_T_11 = fm_div_t2 * fm_col; // @[control.scala 582:56]
  wire [18:0] _ifm_send_len_T_12 = {_ifm_send_len_T_11, 3'h0}; // @[control.scala 582:66]
  wire [18:0] _GEN_30 = _T_17 ? _ifm_send_len_T_6 : _ifm_send_len_T_12; // @[control.scala 576:58 578:42 582:42]
  wire [5:0] _GEN_31 = _T_17 ? fm_div_t1 : fm_div_t2; // @[control.scala 576:58 579:58 583:58]
  wire [18:0] _GEN_33 = _T_16 ? _ifm_send_len_T_2 : _GEN_30; // @[control.scala 572:54 574:42]
  wire [5:0] _GEN_34 = _T_16 ? fm_res_t1 : _GEN_31; // @[control.scala 572:54 575:58]
  wire [15:0] _ifm_send_len_T_13 = fm_res * fm_col; // @[control.scala 588:53]
  wire [18:0] _ifm_send_len_T_14 = {_ifm_send_len_T_13, 3'h0}; // @[control.scala 588:63]
  wire [31:0] _GEN_35 = _T_16 ? fm_row_fm_resxfm_col : iter_div_prexfm_div_col; // @[control.scala 586:54 587:45 591:45]
  wire [18:0] _GEN_36 = _T_16 ? _ifm_send_len_T_14 : _ifm_send_len_T_4; // @[control.scala 586:54 588:42 592:42]
  wire [5:0] _GEN_37 = _T_16 ? fm_res : fm_div; // @[control.scala 586:54 589:59 593:59]
  wire [31:0] _GEN_38 = p_is_1 ? _GEN_22 : _GEN_35; // @[control.scala 571:35]
  wire [18:0] _GEN_39 = p_is_1 ? _GEN_33 : _GEN_36; // @[control.scala 571:35]
  wire [5:0] _GEN_40 = p_is_1 ? _GEN_34 : _GEN_37; // @[control.scala 571:35]
  wire [31:0] _GEN_41 = current_layer_is_conv ? _GEN_25 : _GEN_38; // @[control.scala 553:29]
  wire [31:0] _GEN_42 = current_layer_is_conv ? _GEN_26 : {{13'd0}, _GEN_39}; // @[control.scala 553:29]
  wire [7:0] _GEN_43 = current_layer_is_conv ? _GEN_27 : {{2'd0}, _GEN_40}; // @[control.scala 553:29]
  wire [31:0] _GEN_44 = current_layer_is_conv ? _GEN_28 : reg_linebuffer_sel; // @[control.scala 553:29 596:32]
  wire [31:0] _GEN_45 = fm_div_cnt == 8'h1 ? 32'h0 : _GEN_41; // @[control.scala 543:38 545:33]
  wire [31:0] _GEN_46 = fm_div_cnt == 8'h1 ? {{10'd0}, _ifm_send_len_T} : _GEN_42; // @[control.scala 543:38 548:30]
  wire [9:0] _GEN_47 = fm_div_cnt == 8'h1 ? fm_col : {{2'd0}, _GEN_43}; // @[control.scala 543:38 550:47]
  wire [31:0] _GEN_48 = fm_div_cnt == 8'h1 ? reg_static : _GEN_44; // @[control.scala 161:29 543:38]
  wire [31:0] _reg_static_T_1 = reg_static | 32'h40; // @[control.scala 606:46]
  wire [31:0] _reg_static_T_2 = _reg_static_T_1 | 32'h80; // @[control.scala 606:59]
  wire [31:0] _GEN_49 = ifm_batch == 13'h1 ? _reg_static_T_2 : _reg_static_T_1; // @[control.scala 605:40 606:32 608:32]
  wire [12:0] _T_25 = ifm_batch - 13'h1; // @[control.scala 610:52]
  wire  _T_26 = iter_ifm_post == _T_25; // @[control.scala 610:38]
  wire [31:0] _reg_static_T_4 = reg_static | 32'h80; // @[control.scala 611:42]
  wire [31:0] _GEN_50 = iter_ifm_post == _T_25 ? _reg_static_T_4 : reg_static; // @[control.scala 610:59 611:28 161:29]
  wire [31:0] _GEN_51 = iter_ifm_post == 13'h0 ? _GEN_49 : _GEN_50; // @[control.scala 604:41]
  wire  _T_28 = ~last_buf_sel; // @[control.scala 616:18]
  wire [31:0] _reg_static_T_5 = reg_static | 32'h100; // @[control.scala 617:42]
  wire [31:0] _GEN_52 = ~last_buf_sel ? _reg_static_T_5 : reg_static; // @[control.scala 616:33 617:28 161:29]
  wire [31:0] _reg_static_T_6 = reg_static | 32'h10000; // @[control.scala 624:42]
  wire [31:0] _reg_static_T_7 = _reg_static_T_6 | 32'h20000; // @[control.scala 624:60]
  wire [31:0] _reg_static_T_9 = reg_static | 32'h20000; // @[control.scala 628:42]
  wire [31:0] _GEN_53 = skip_act ? _reg_static_T_9 : reg_static; // @[control.scala 627:34 628:28 161:29]
  wire [31:0] _GEN_54 = upsample_en ? _reg_static_T_6 : _GEN_53; // @[control.scala 625:37 626:28]
  wire [31:0] _GEN_55 = upsample_en & skip_act ? _reg_static_T_7 : _GEN_54; // @[control.scala 623:43 624:28]
  wire [31:0] _reg_static_T_12 = {the_number_of_row_transferred,reg_static[23:16],3'h7,reg_static[12:0]}; // @[Cat.scala 33:92]
  wire [31:0] _reg_static_T_14 = {the_number_of_row_transferred,reg_static[23:0]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_56 = p_is_1 ? _reg_static_T_12 : _reg_static_T_14; // @[control.scala 634:31 635:32 637:32]
  wire [31:0] _reg_static_T_17 = {the_number_of_row_transferred,reg_static[23:16],3'h5,reg_static[12:0]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_57 = p_is_1 ? _reg_static_T_17 : _reg_static_T_14; // @[control.scala 641:35 642:36 644:36]
  wire  _T_34 = _iter_div_post_t_T_1 == 13'h1; // @[control.scala 646:44]
  wire [31:0] _reg_static_T_22 = {the_number_of_row_transferred,reg_static[23:16],3'h6,reg_static[12:0]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_58 = p_is_1 ? _reg_static_T_22 : _reg_static_T_14; // @[control.scala 647:35 648:36 650:36]
  wire [31:0] _reg_static_T_27 = {the_number_of_row_transferred,reg_static[23:16],3'h4,reg_static[12:0]}; // @[Cat.scala 33:92]
  wire [31:0] _GEN_59 = p_is_1 ? _reg_static_T_27 : _reg_static_T_14; // @[control.scala 653:35 654:36 656:36]
  wire [31:0] _GEN_60 = _iter_div_post_t_T_1 == 13'h1 ? _GEN_58 : _GEN_59; // @[control.scala 646:53]
  wire [31:0] _GEN_61 = iter_div_post == 13'h0 ? _GEN_57 : _GEN_60; // @[control.scala 640:45]
  wire [31:0] _GEN_62 = _T_15 ? _GEN_56 : _GEN_61; // @[control.scala 633:38]
  wire  _T_39 = iter_ofm_post_t == 13'h1 & _T_34 & _ofm_write_disable_T; // @[control.scala 661:69]
  wire [19:0] _GEN_63 = bottleneck_ready ? 20'h80200 : 20'h210; // @[control.scala 662:39 663:30 665:30]
  wire  _T_44 = iter_ofm_pre == 13'h0 & _T_17 & iter_ifm_pre == 13'h0; // @[control.scala 667:69]
  wire [19:0] _GEN_64 = bottleneck_ready ? 20'h80201 : 20'h211; // @[control.scala 670:39 671:30 673:30]
  wire [19:0] _GEN_65 = iter_ofm_pre == 13'h0 & _T_17 & iter_ifm_pre == 13'h0 ? 20'h201 : _GEN_64; // @[control.scala 667:94 668:26]
  wire [19:0] _GEN_66 = iter_ofm_post_t == 13'h1 & _T_34 & _ofm_write_disable_T ? _GEN_63 : _GEN_65; // @[control.scala 661:97]
  wire [31:0] _GEN_67 = ifm_send_task_enable ? ifm_addr_send : reg_t_4; // @[control.scala 684:40 685:26 160:37]
  wire [31:0] _GEN_68 = ifm_send_task_enable ? ifm_send_len : reg_t_5; // @[control.scala 684:40 686:26 160:37]
  wire [31:0] _reg_t_3_T_2 = {bia_addr_read,weight_sel,wgt_addr_read[12:0]}; // @[Cat.scala 33:92]
  wire [31:0] _reg_t_0_T_4 = reg_static | reg_task; // @[control.scala 690:36]
  wire [5:0] _GEN_70 = cnt_t_is_5 ? 6'hf : state; // @[control.scala 695:30 697:23 436:24]
  wire [31:0] _GEN_71 = cnt_t_is_5 ? reg_static : reg_t_0; // @[control.scala 695:30 698:26 160:37]
  wire  _GEN_72 = bottleneck_transfer ? 1'h0 : bottleneck_transfer; // @[control.scala 295:38 707:43 708:41]
  wire  _GEN_73 = bottleneck_transfer | bottleneck_ready; // @[control.scala 296:35 707:43 709:38]
  wire  _GEN_74 = bottleneck_ready ? 1'h0 : _GEN_73; // @[control.scala 711:40 712:38]
  wire [4:0] _GEN_75 = ap_done_up ? 5'h10 : 5'hf; // @[control.scala 705:30 706:23 715:23]
  wire  _GEN_76 = ap_done_up ? _GEN_72 : bottleneck_transfer; // @[control.scala 705:30 295:38]
  wire  _GEN_77 = ap_done_up ? _GEN_74 : bottleneck_ready; // @[control.scala 705:30 296:35]
  wire  _T_58 = ~first_ofm_recv_stop & _ofm_write_disable_T & _ofm_write_disable_T_1 & (~_skip_act_T_3 | _skip_act_T_3
     & _T_34); // @[control.scala 721:91]
  wire [4:0] _GEN_79 = ~first_ofm_recv_stop & _ofm_write_disable_T & _ofm_write_disable_T_1 & (~_skip_act_T_3 |
    _skip_act_T_3 & _T_34) ? 5'h11 : 5'h13; // @[control.scala 721:156 725:23 728:23]
  wire  _GEN_80 = ~first_ofm_recv_stop & _ofm_write_disable_T & _ofm_write_disable_T_1 & (~_skip_act_T_3 | _skip_act_T_3
     & _T_34) & first_ofm_recv_stop; // @[control.scala 721:156 422:38 729:37]
  wire [31:0] _ofm_addr_fmbase_T = iter_ofm_post * fm_size_output; // @[control.scala 733:46]
  wire [21:0] _ofm_recv_len_T = {fm_size_output, 3'h0}; // @[control.scala 737:47]
  wire [31:0] _GEN_81 = _T_15 ? 32'h0 : ofm_addr_offset; // @[control.scala 735:36 736:33 366:34]
  wire [31:0] _GEN_82 = _T_15 ? {{10'd0}, _ofm_recv_len_T} : ofm_recv_len; // @[control.scala 735:36 737:30 367:31]
  wire [4:0] _GEN_83 = _T_15 ? 5'h13 : 5'h12; // @[control.scala 735:36 738:23 740:23]
  wire [15:0] _ofm_recv_len_T_1 = fm_res_output * fm_col_output; // @[control.scala 747:48]
  wire [18:0] _ofm_recv_len_T_2 = {_ofm_recv_len_T_1, 3'h0}; // @[control.scala 747:65]
  wire [15:0] _ofm_recv_len_T_3 = fm_div_output * fm_col_output; // @[control.scala 750:48]
  wire [18:0] _ofm_recv_len_T_4 = {_ofm_recv_len_T_3, 3'h0}; // @[control.scala 750:65]
  wire [31:0] _GEN_84 = _T_34 ? fm_row_res_outputxfm_col_output : iter_div_postxfm_col_output; // @[control.scala 745:43 746:33 749:33]
  wire [18:0] _GEN_85 = _T_34 ? _ofm_recv_len_T_2 : _ofm_recv_len_T_4; // @[control.scala 745:43 747:30 750:30]
  wire  _T_67 = wgt_ddr_read_en & _T_34 & _T_9; // @[control.scala 756:61]
  wire [31:0] _GEN_2846 = {{12'd0}, _reg_t_5_T_6}; // @[control.scala 758:48]
  wire [31:0] _wgt_addr_send_T_7 = wgt_addr_send + _GEN_2846; // @[control.scala 758:48]
  wire [31:0] _GEN_87 = wgt_ddr_read_en & _T_34 & _T_9 ? _wgt_addr_send_T_7 : wgt_addr_send; // @[control.scala 756:89 758:31 178:32]
  wire [15:0] _GEN_88 = wgt_ddr_read_en & _T_34 & _T_9 ? 16'h0 : wgt_addr_read; // @[control.scala 756:89 759:31 179:32]
  wire [5:0] _GEN_89 = ~ofm_recv_task_enable ? 6'h14 : 6'h20; // @[control.scala 764:41 765:23 767:23]
  wire [12:0] _iter_ifm_pre_T_1 = iter_ifm_pre + 13'h1; // @[control.scala 777:46]
  wire [4:0] _GEN_90 = bottleneck_transfer ? 5'h19 : 5'h15; // @[control.scala 774:38 775:23 778:23]
  wire [12:0] _GEN_91 = bottleneck_transfer ? iter_ifm_pre : _iter_ifm_pre_T_1; // @[control.scala 192:31 774:38 777:30]
  wire  _bottleneck_transfer_T_1 = bottleneck_en & iter_ifm_pre_t == 13'h1; // @[control.scala 783:50]
  wire  _T_71 = iter_ifm_pre == ifm_batch; // @[control.scala 784:31]
  wire [12:0] _iter_div_pre_T_1 = iter_div_pre + 13'h1; // @[control.scala 786:46]
  wire [12:0] _GEN_92 = iter_ifm_pre == ifm_batch ? 13'h0 : iter_ifm_pre; // @[control.scala 784:46 785:30 192:31]
  wire [12:0] _GEN_93 = iter_ifm_pre == ifm_batch ? _iter_div_pre_T_1 : iter_div_pre; // @[control.scala 784:46 786:30 195:31]
  wire [4:0] _GEN_94 = iter_ifm_pre == ifm_batch ? 5'h16 : 5'h17; // @[control.scala 784:46 787:23 789:23]
  wire [12:0] _iter_ofm_pre_T_1 = iter_ofm_pre + 13'h1; // @[control.scala 795:46]
  wire [12:0] _GEN_95 = iter_div_pre == _GEN_2833 ? 13'h0 : iter_div_pre; // @[control.scala 793:47 794:30 195:31]
  wire [12:0] _GEN_96 = iter_div_pre == _GEN_2833 ? _iter_ofm_pre_T_1 : iter_ofm_pre; // @[control.scala 793:47 795:30 194:31]
  wire [4:0] _GEN_98 = _T_13 ? 5'h18 : 5'h1a; // @[control.scala 801:97 803:23 806:23]
  wire [31:0] _GEN_131 = _T_15 ? 32'h0 : _GEN_84; // @[control.scala 868:38 869:33]
  wire [21:0] _GEN_132 = _T_15 ? _ofm_recv_len_T : {{3'd0}, _GEN_85}; // @[control.scala 868:38 870:30]
  wire [9:0] _GEN_147 = _T_44 ? 10'h201 : 10'h211; // @[control.scala 945:94 946:26 948:26]
  wire [9:0] _GEN_148 = _T_39 ? 10'h210 : _GEN_147; // @[control.scala 943:97 944:26]
  wire [25:0] _wgt_addr_read_t_T_1 = iter_ofm_post * ifm_batch; // @[control.scala 959:54]
  wire [25:0] _GEN_2850 = {{13'd0}, iter_ifm_post}; // @[control.scala 959:66]
  wire [25:0] _wgt_addr_read_t_T_3 = _wgt_addr_read_t_T_1 + _GEN_2850; // @[control.scala 959:66]
  wire [25:0] _GEN_149 = ifm_batch_is_exactly_divided_by_WEIGHT_LEN ? _wgt_addr_read_t_T_3 : {{13'd0}, iter_ifm_post}; // @[control.scala 958:65 959:37 961:37]
  wire [25:0] _GEN_150 = k_is_1 ? {{16'd0}, iter_ifm_post[12:3]} : _GEN_149; // @[control.scala 954:25 955:32]
  wire [2:0] _GEN_151 = k_is_1 ? iter_ifm_post[2:0] : weight_sel; // @[control.scala 954:25 274:27 956:27]
  wire [15:0] _wgt_addr_read_T = wgt_addr_read_t & 16'h7f; // @[control.scala 967:46]
  wire [7:0] _wgt_ddr_read_en_T_4 = weight_len - 8'h1; // @[control.scala 969:103]
  wire [15:0] _GEN_2851 = {{8'd0}, _wgt_ddr_read_en_T_4}; // @[control.scala 969:87]
  wire  _wgt_ddr_read_en_T_6 = k_is_1 ? _T_26 : wgt_addr_read == _GEN_2851; // @[control.scala 969:33]
  wire [5:0] _GEN_152 = ~pool_en ? 6'h23 : 6'h21; // @[control.scala 976:31 977:27 979:27]
  wire [5:0] _GEN_153 = ofm_recv_task_enable ? _GEN_152 : 6'h32; // @[control.scala 975:40 983:23]
  wire [31:0] _reg_t_0_T_5 = reg_t_0 | 32'h20; // @[control.scala 987:34]
  wire [5:0] _GEN_154 = io_pool_finish_edge ? 6'h23 : 6'h22; // @[control.scala 991:30 992:22 994:23]
  wire [31:0] _reg_t_0_T_6 = reg_static | 32'h2; // @[control.scala 1005:36]
  wire [31:0] _reg_t_0_T_7 = _reg_t_0_T_6 | 32'h200; // @[control.scala 1005:50]
  wire [5:0] _GEN_156 = cnt_t_is_5 ? 6'h25 : state; // @[control.scala 1010:30 1013:23 436:24]
  wire [2:0] _GEN_2852 = {{1'd0}, pool_cnt}; // @[control.scala 1026:34]
  wire [1:0] _pool_cnt_T_1 = pool_cnt + 2'h1; // @[control.scala 1030:43]
  wire [1:0] _GEN_157 = _GEN_2852 == 3'h4 ? 2'h0 : _pool_cnt_T_1; // @[control.scala 1026:69 1027:33 1030:33]
  wire [5:0] _GEN_158 = _GEN_2852 == 3'h4 ? 6'h26 : 6'h23; // @[control.scala 1026:69 1028:31 1031:30]
  wire [1:0] _GEN_159 = pool_en ? _GEN_157 : pool_cnt; // @[control.scala 1023:30 290:27]
  wire [5:0] _GEN_160 = pool_en ? _GEN_158 : 6'h26; // @[control.scala 1023:30 1034:27]
  wire [1:0] _GEN_161 = ap_done_up ? _GEN_159 : pool_cnt; // @[control.scala 1022:30 290:27]
  wire [5:0] _GEN_162 = ap_done_up ? _GEN_160 : 6'h25; // @[control.scala 1022:30 1037:23]
  wire [5:0] _GEN_163 = bottleneck_transfer ? 6'h2b : 6'h27; // @[control.scala 1049:42 1050:27 1053:27]
  wire [5:0] _GEN_165 = _T_39 ? 6'h36 : _GEN_163; // @[control.scala 1042:97 1043:23]
  wire [12:0] _GEN_166 = _T_39 ? iter_ifm_post : iter_ifm_pre; // @[control.scala 1042:97 1045:31 196:32]
  wire [12:0] _GEN_167 = _T_39 ? iter_div_post : iter_div_pre; // @[control.scala 1042:97 1046:31 198:32]
  wire [12:0] _GEN_168 = _T_39 ? iter_ofm_post : iter_ofm_pre; // @[control.scala 1042:97 1047:31 197:32]
  wire [12:0] _GEN_169 = _T_39 ? iter_ifm_pre : _GEN_91; // @[control.scala 1042:97 192:31]
  wire [5:0] _GEN_172 = _T_71 ? 6'h28 : 6'h29; // @[control.scala 1060:46 1063:23 1065:23]
  wire [5:0] _GEN_176 = _T_13 ? 6'h2a : 6'h2c; // @[control.scala 1076:97 1078:23 1081:23]
  wire [5:0] _GEN_230 = wgt_send_task_enable ? 6'h33 : 6'hd; // @[control.scala 1246:40 1247:23 1249:23]
  wire [5:0] _GEN_232 = cnt_t_is_5 ? 6'h35 : state; // @[control.scala 1260:30 1262:23 436:24]
  wire [5:0] _GEN_233 = ap_done_up ? 6'hd : 6'h35; // @[control.scala 1269:30 1270:23 1272:23]
  wire  _GEN_234 = current_layer == 5'h16 ? ~ifm_sel : ifm_sel; // @[control.scala 1280:56 1281:25 379:24]
  wire  _GEN_236 = current_layer == 5'h16 ? ~resize_load_t : resize_load_t; // @[control.scala 1280:56 1286:31 420:32]
  wire  _GEN_237 = current_layer == 5'h16 | yolo_finish; // @[control.scala 1280:56 1288:29 40:28]
  wire  _GEN_238 = 6'h36 == state ? _GEN_234 : ifm_sel; // @[control.scala 438:19 379:24]
  wire [5:0] _GEN_239 = 6'h36 == state ? 6'h0 : state; // @[control.scala 438:19 1294:23 436:24]
  wire  _GEN_240 = 6'h36 == state ? _GEN_236 : resize_load_t; // @[control.scala 438:19 420:32]
  wire  _GEN_241 = 6'h36 == state ? _GEN_237 : yolo_finish; // @[control.scala 438:19 40:28]
  wire  _GEN_242 = 6'h36 == state | conv_finish; // @[control.scala 438:19 1292:29 71:30]
  wire [5:0] _GEN_243 = 6'h35 == state ? _GEN_233 : _GEN_239; // @[control.scala 438:19]
  wire  _GEN_244 = 6'h35 == state ? ifm_sel : _GEN_238; // @[control.scala 438:19 379:24]
  wire  _GEN_245 = 6'h35 == state ? resize_load_t : _GEN_240; // @[control.scala 438:19 420:32]
  wire  _GEN_246 = 6'h35 == state ? yolo_finish : _GEN_241; // @[control.scala 438:19 40:28]
  wire  _GEN_247 = 6'h35 == state ? conv_finish : _GEN_242; // @[control.scala 438:19 71:30]
  wire [4:0] _GEN_248 = 6'h34 == state ? _GEN_2 : cnt_t; // @[control.scala 438:19 163:24]
  wire [5:0] _GEN_249 = 6'h34 == state ? _GEN_232 : _GEN_243; // @[control.scala 438:19]
  wire [31:0] _GEN_250 = 6'h34 == state ? _GEN_11 : reg_t_0; // @[control.scala 438:19 160:37]
  wire  _GEN_251 = 6'h34 == state ? ifm_sel : _GEN_244; // @[control.scala 438:19 379:24]
  wire  _GEN_252 = 6'h34 == state ? resize_load_t : _GEN_245; // @[control.scala 438:19 420:32]
  wire  _GEN_253 = 6'h34 == state ? yolo_finish : _GEN_246; // @[control.scala 438:19 40:28]
  wire  _GEN_254 = 6'h34 == state ? conv_finish : _GEN_247; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_255 = 6'h33 == state ? wgt_addr_send : reg_t_4; // @[control.scala 438:19 1253:22 160:37]
  wire [31:0] _GEN_256 = 6'h33 == state ? {{12'd0}, _reg_t_5_T_6} : reg_t_5; // @[control.scala 438:19 1254:22 160:37]
  wire [31:0] _GEN_257 = 6'h33 == state ? 32'h205 : _GEN_250; // @[control.scala 438:19 1255:22]
  wire [4:0] _GEN_258 = 6'h33 == state ? 5'h0 : _GEN_248; // @[control.scala 1256:19 438:19]
  wire [5:0] _GEN_259 = 6'h33 == state ? 6'h34 : _GEN_249; // @[control.scala 1257:19 438:19]
  wire  _GEN_260 = 6'h33 == state ? ifm_sel : _GEN_251; // @[control.scala 438:19 379:24]
  wire  _GEN_261 = 6'h33 == state ? resize_load_t : _GEN_252; // @[control.scala 438:19 420:32]
  wire  _GEN_262 = 6'h33 == state ? yolo_finish : _GEN_253; // @[control.scala 438:19 40:28]
  wire  _GEN_263 = 6'h33 == state ? conv_finish : _GEN_254; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_264 = 6'h32 == state ? _GEN_230 : _GEN_259; // @[control.scala 438:19]
  wire [31:0] _GEN_265 = 6'h32 == state ? reg_t_4 : _GEN_255; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_266 = 6'h32 == state ? reg_t_5 : _GEN_256; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_267 = 6'h32 == state ? reg_t_0 : _GEN_257; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_268 = 6'h32 == state ? cnt_t : _GEN_258; // @[control.scala 438:19 163:24]
  wire  _GEN_269 = 6'h32 == state ? ifm_sel : _GEN_260; // @[control.scala 438:19 379:24]
  wire  _GEN_270 = 6'h32 == state ? resize_load_t : _GEN_261; // @[control.scala 438:19 420:32]
  wire  _GEN_271 = 6'h32 == state ? yolo_finish : _GEN_262; // @[control.scala 438:19 40:28]
  wire  _GEN_272 = 6'h32 == state ? conv_finish : _GEN_263; // @[control.scala 438:19 71:30]
  wire [15:0] _GEN_273 = 6'h31 == state ? _wgt_addr_read_T : wgt_addr_read; // @[control.scala 438:19 1240:27 179:32]
  wire [15:0] _GEN_274 = 6'h31 == state ? {{3'd0}, iter_ofm_post} : bia_addr_read; // @[control.scala 438:19 1241:27 181:32]
  wire  _GEN_275 = 6'h31 == state ? _wgt_ddr_read_en_T_6 : wgt_ddr_read_en; // @[control.scala 438:19 1242:28 424:32]
  wire [5:0] _GEN_276 = 6'h31 == state ? 6'h32 : _GEN_264; // @[control.scala 1243:19 438:19]
  wire [31:0] _GEN_277 = 6'h31 == state ? reg_t_4 : _GEN_265; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_278 = 6'h31 == state ? reg_t_5 : _GEN_266; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_279 = 6'h31 == state ? reg_t_0 : _GEN_267; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_280 = 6'h31 == state ? cnt_t : _GEN_268; // @[control.scala 438:19 163:24]
  wire  _GEN_281 = 6'h31 == state ? ifm_sel : _GEN_269; // @[control.scala 438:19 379:24]
  wire  _GEN_282 = 6'h31 == state ? resize_load_t : _GEN_270; // @[control.scala 438:19 420:32]
  wire  _GEN_283 = 6'h31 == state ? yolo_finish : _GEN_271; // @[control.scala 438:19 40:28]
  wire  _GEN_284 = 6'h31 == state ? conv_finish : _GEN_272; // @[control.scala 438:19 71:30]
  wire [25:0] _GEN_285 = 6'h30 == state ? _GEN_150 : {{10'd0}, wgt_addr_read_t}; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_286 = 6'h30 == state ? _GEN_151 : weight_sel; // @[control.scala 438:19 274:27]
  wire [5:0] _GEN_287 = 6'h30 == state ? 6'h31 : _GEN_276; // @[control.scala 1237:19 438:19]
  wire [15:0] _GEN_288 = 6'h30 == state ? wgt_addr_read : _GEN_273; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_289 = 6'h30 == state ? bia_addr_read : _GEN_274; // @[control.scala 438:19 181:32]
  wire  _GEN_290 = 6'h30 == state ? wgt_ddr_read_en : _GEN_275; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_291 = 6'h30 == state ? reg_t_4 : _GEN_277; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_292 = 6'h30 == state ? reg_t_5 : _GEN_278; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_293 = 6'h30 == state ? reg_t_0 : _GEN_279; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_294 = 6'h30 == state ? cnt_t : _GEN_280; // @[control.scala 438:19 163:24]
  wire  _GEN_295 = 6'h30 == state ? ifm_sel : _GEN_281; // @[control.scala 438:19 379:24]
  wire  _GEN_296 = 6'h30 == state ? resize_load_t : _GEN_282; // @[control.scala 438:19 420:32]
  wire  _GEN_297 = 6'h30 == state ? yolo_finish : _GEN_283; // @[control.scala 438:19 40:28]
  wire  _GEN_298 = 6'h30 == state ? conv_finish : _GEN_284; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_299 = 6'h2f == state ? _GEN_62 : reg_static; // @[control.scala 438:19 161:29]
  wire [31:0] _GEN_300 = 6'h2f == state ? {{22'd0}, _GEN_148} : reg_task; // @[control.scala 438:19 162:27]
  wire [5:0] _GEN_301 = 6'h2f == state ? 6'h30 : _GEN_287; // @[control.scala 1224:19 438:19]
  wire [25:0] _GEN_302 = 6'h2f == state ? {{10'd0}, wgt_addr_read_t} : _GEN_285; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_303 = 6'h2f == state ? weight_sel : _GEN_286; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_304 = 6'h2f == state ? wgt_addr_read : _GEN_288; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_305 = 6'h2f == state ? bia_addr_read : _GEN_289; // @[control.scala 438:19 181:32]
  wire  _GEN_306 = 6'h2f == state ? wgt_ddr_read_en : _GEN_290; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_307 = 6'h2f == state ? reg_t_4 : _GEN_291; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_308 = 6'h2f == state ? reg_t_5 : _GEN_292; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_309 = 6'h2f == state ? reg_t_0 : _GEN_293; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_310 = 6'h2f == state ? cnt_t : _GEN_294; // @[control.scala 438:19 163:24]
  wire  _GEN_311 = 6'h2f == state ? ifm_sel : _GEN_295; // @[control.scala 438:19 379:24]
  wire  _GEN_312 = 6'h2f == state ? resize_load_t : _GEN_296; // @[control.scala 438:19 420:32]
  wire  _GEN_313 = 6'h2f == state ? yolo_finish : _GEN_297; // @[control.scala 438:19 40:28]
  wire  _GEN_314 = 6'h2f == state ? conv_finish : _GEN_298; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_315 = 6'h2e == state ? _GEN_55 : _GEN_299; // @[control.scala 438:19]
  wire [5:0] _GEN_316 = 6'h2e == state ? 6'h2f : _GEN_301; // @[control.scala 1187:18 438:19]
  wire [31:0] _GEN_317 = 6'h2e == state ? reg_task : _GEN_300; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_318 = 6'h2e == state ? {{10'd0}, wgt_addr_read_t} : _GEN_302; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_319 = 6'h2e == state ? weight_sel : _GEN_303; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_320 = 6'h2e == state ? wgt_addr_read : _GEN_304; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_321 = 6'h2e == state ? bia_addr_read : _GEN_305; // @[control.scala 438:19 181:32]
  wire  _GEN_322 = 6'h2e == state ? wgt_ddr_read_en : _GEN_306; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_323 = 6'h2e == state ? reg_t_4 : _GEN_307; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_324 = 6'h2e == state ? reg_t_5 : _GEN_308; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_325 = 6'h2e == state ? reg_t_0 : _GEN_309; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_326 = 6'h2e == state ? cnt_t : _GEN_310; // @[control.scala 438:19 163:24]
  wire  _GEN_327 = 6'h2e == state ? ifm_sel : _GEN_311; // @[control.scala 438:19 379:24]
  wire  _GEN_328 = 6'h2e == state ? resize_load_t : _GEN_312; // @[control.scala 438:19 420:32]
  wire  _GEN_329 = 6'h2e == state ? yolo_finish : _GEN_313; // @[control.scala 438:19 40:28]
  wire  _GEN_330 = 6'h2e == state ? conv_finish : _GEN_314; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_331 = 6'h2d == state ? _GEN_52 : _GEN_315; // @[control.scala 438:19]
  wire  _GEN_332 = 6'h2d == state ? _T_28 : last_buf_sel; // @[control.scala 438:19 1176:26 182:31]
  wire [5:0] _GEN_333 = 6'h2d == state ? 6'h2e : _GEN_316; // @[control.scala 1177:19 438:19]
  wire [31:0] _GEN_334 = 6'h2d == state ? reg_task : _GEN_317; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_335 = 6'h2d == state ? {{10'd0}, wgt_addr_read_t} : _GEN_318; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_336 = 6'h2d == state ? weight_sel : _GEN_319; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_337 = 6'h2d == state ? wgt_addr_read : _GEN_320; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_338 = 6'h2d == state ? bia_addr_read : _GEN_321; // @[control.scala 438:19 181:32]
  wire  _GEN_339 = 6'h2d == state ? wgt_ddr_read_en : _GEN_322; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_340 = 6'h2d == state ? reg_t_4 : _GEN_323; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_341 = 6'h2d == state ? reg_t_5 : _GEN_324; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_342 = 6'h2d == state ? reg_t_0 : _GEN_325; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_343 = 6'h2d == state ? cnt_t : _GEN_326; // @[control.scala 438:19 163:24]
  wire  _GEN_344 = 6'h2d == state ? ifm_sel : _GEN_327; // @[control.scala 438:19 379:24]
  wire  _GEN_345 = 6'h2d == state ? resize_load_t : _GEN_328; // @[control.scala 438:19 420:32]
  wire  _GEN_346 = 6'h2d == state ? yolo_finish : _GEN_329; // @[control.scala 438:19 40:28]
  wire  _GEN_347 = 6'h2d == state ? conv_finish : _GEN_330; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_348 = 6'h2c == state ? _GEN_51 : _GEN_331; // @[control.scala 438:19]
  wire [5:0] _GEN_349 = 6'h2c == state ? 6'h2d : _GEN_333; // @[control.scala 1169:19 438:19]
  wire  _GEN_350 = 6'h2c == state ? last_buf_sel : _GEN_332; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_351 = 6'h2c == state ? reg_task : _GEN_334; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_352 = 6'h2c == state ? {{10'd0}, wgt_addr_read_t} : _GEN_335; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_353 = 6'h2c == state ? weight_sel : _GEN_336; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_354 = 6'h2c == state ? wgt_addr_read : _GEN_337; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_355 = 6'h2c == state ? bia_addr_read : _GEN_338; // @[control.scala 438:19 181:32]
  wire  _GEN_356 = 6'h2c == state ? wgt_ddr_read_en : _GEN_339; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_357 = 6'h2c == state ? reg_t_4 : _GEN_340; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_358 = 6'h2c == state ? reg_t_5 : _GEN_341; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_359 = 6'h2c == state ? reg_t_0 : _GEN_342; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_360 = 6'h2c == state ? cnt_t : _GEN_343; // @[control.scala 438:19 163:24]
  wire  _GEN_361 = 6'h2c == state ? ifm_sel : _GEN_344; // @[control.scala 438:19 379:24]
  wire  _GEN_362 = 6'h2c == state ? resize_load_t : _GEN_345; // @[control.scala 438:19 420:32]
  wire  _GEN_363 = 6'h2c == state ? yolo_finish : _GEN_346; // @[control.scala 438:19 40:28]
  wire  _GEN_364 = 6'h2c == state ? conv_finish : _GEN_347; // @[control.scala 438:19 71:30]
  wire  _GEN_365 = 6'h2b == state | ifm_send_task_enable; // @[control.scala 438:19 1142:34 357:39]
  wire [31:0] _GEN_366 = 6'h2b == state ? _ofm_addr_fmbase_T : ifm_addr_fmbase; // @[control.scala 438:19 1143:29 362:34]
  wire [31:0] _GEN_367 = 6'h2b == state ? _GEN_131 : ifm_addr_offset; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_368 = 6'h2b == state ? {{10'd0}, _GEN_132} : ifm_send_len; // @[control.scala 438:19 364:31]
  wire [5:0] _GEN_369 = 6'h2b == state ? 6'h2c : _GEN_349; // @[control.scala 1156:19 438:19]
  wire [31:0] _GEN_370 = 6'h2b == state ? reg_static : _GEN_348; // @[control.scala 438:19 161:29]
  wire  _GEN_371 = 6'h2b == state ? last_buf_sel : _GEN_350; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_372 = 6'h2b == state ? reg_task : _GEN_351; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_373 = 6'h2b == state ? {{10'd0}, wgt_addr_read_t} : _GEN_352; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_374 = 6'h2b == state ? weight_sel : _GEN_353; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_375 = 6'h2b == state ? wgt_addr_read : _GEN_354; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_376 = 6'h2b == state ? bia_addr_read : _GEN_355; // @[control.scala 438:19 181:32]
  wire  _GEN_377 = 6'h2b == state ? wgt_ddr_read_en : _GEN_356; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_378 = 6'h2b == state ? reg_t_4 : _GEN_357; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_379 = 6'h2b == state ? reg_t_5 : _GEN_358; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_380 = 6'h2b == state ? reg_t_0 : _GEN_359; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_381 = 6'h2b == state ? cnt_t : _GEN_360; // @[control.scala 438:19 163:24]
  wire  _GEN_382 = 6'h2b == state ? ifm_sel : _GEN_361; // @[control.scala 438:19 379:24]
  wire  _GEN_383 = 6'h2b == state ? resize_load_t : _GEN_362; // @[control.scala 438:19 420:32]
  wire  _GEN_384 = 6'h2b == state ? yolo_finish : _GEN_363; // @[control.scala 438:19 40:28]
  wire  _GEN_385 = 6'h2b == state ? conv_finish : _GEN_364; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_386 = 6'h2a == state ? _ifm_addr_fmbase_T : _GEN_366; // @[control.scala 438:19 1086:29]
  wire [31:0] _GEN_387 = 6'h2a == state ? _GEN_45 : _GEN_367; // @[control.scala 438:19]
  wire [31:0] _GEN_388 = 6'h2a == state ? _GEN_46 : _GEN_368; // @[control.scala 438:19]
  wire [9:0] _GEN_389 = 6'h2a == state ? _GEN_47 : {{2'd0}, the_number_of_row_transferred}; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_390 = 6'h2a == state ? _GEN_48 : _GEN_370; // @[control.scala 438:19]
  wire [5:0] _GEN_391 = 6'h2a == state ? 6'h2c : _GEN_369; // @[control.scala 1139:19 438:19]
  wire  _GEN_392 = 6'h2a == state ? ifm_send_task_enable : _GEN_365; // @[control.scala 438:19 357:39]
  wire  _GEN_393 = 6'h2a == state ? last_buf_sel : _GEN_371; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_394 = 6'h2a == state ? reg_task : _GEN_372; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_395 = 6'h2a == state ? {{10'd0}, wgt_addr_read_t} : _GEN_373; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_396 = 6'h2a == state ? weight_sel : _GEN_374; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_397 = 6'h2a == state ? wgt_addr_read : _GEN_375; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_398 = 6'h2a == state ? bia_addr_read : _GEN_376; // @[control.scala 438:19 181:32]
  wire  _GEN_399 = 6'h2a == state ? wgt_ddr_read_en : _GEN_377; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_400 = 6'h2a == state ? reg_t_4 : _GEN_378; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_401 = 6'h2a == state ? reg_t_5 : _GEN_379; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_402 = 6'h2a == state ? reg_t_0 : _GEN_380; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_403 = 6'h2a == state ? cnt_t : _GEN_381; // @[control.scala 438:19 163:24]
  wire  _GEN_404 = 6'h2a == state ? ifm_sel : _GEN_382; // @[control.scala 438:19 379:24]
  wire  _GEN_405 = 6'h2a == state ? resize_load_t : _GEN_383; // @[control.scala 438:19 420:32]
  wire  _GEN_406 = 6'h2a == state ? yolo_finish : _GEN_384; // @[control.scala 438:19 40:28]
  wire  _GEN_407 = 6'h2a == state ? conv_finish : _GEN_385; // @[control.scala 438:19 71:30]
  wire  _GEN_408 = 6'h29 == state ? _T_13 : _GEN_392; // @[control.scala 438:19]
  wire [5:0] _GEN_409 = 6'h29 == state ? _GEN_176 : _GEN_391; // @[control.scala 438:19]
  wire [31:0] _GEN_410 = 6'h29 == state ? ifm_addr_fmbase : _GEN_386; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_411 = 6'h29 == state ? ifm_addr_offset : _GEN_387; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_412 = 6'h29 == state ? ifm_send_len : _GEN_388; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_413 = 6'h29 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_389; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_414 = 6'h29 == state ? reg_static : _GEN_390; // @[control.scala 438:19 161:29]
  wire  _GEN_415 = 6'h29 == state ? last_buf_sel : _GEN_393; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_416 = 6'h29 == state ? reg_task : _GEN_394; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_417 = 6'h29 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_395; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_418 = 6'h29 == state ? weight_sel : _GEN_396; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_419 = 6'h29 == state ? wgt_addr_read : _GEN_397; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_420 = 6'h29 == state ? bia_addr_read : _GEN_398; // @[control.scala 438:19 181:32]
  wire  _GEN_421 = 6'h29 == state ? wgt_ddr_read_en : _GEN_399; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_422 = 6'h29 == state ? reg_t_4 : _GEN_400; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_423 = 6'h29 == state ? reg_t_5 : _GEN_401; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_424 = 6'h29 == state ? reg_t_0 : _GEN_402; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_425 = 6'h29 == state ? cnt_t : _GEN_403; // @[control.scala 438:19 163:24]
  wire  _GEN_426 = 6'h29 == state ? ifm_sel : _GEN_404; // @[control.scala 438:19 379:24]
  wire  _GEN_427 = 6'h29 == state ? resize_load_t : _GEN_405; // @[control.scala 438:19 420:32]
  wire  _GEN_428 = 6'h29 == state ? yolo_finish : _GEN_406; // @[control.scala 438:19 40:28]
  wire  _GEN_429 = 6'h29 == state ? conv_finish : _GEN_407; // @[control.scala 438:19 71:30]
  wire [12:0] _GEN_430 = 6'h28 == state ? _GEN_95 : iter_div_pre; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_431 = 6'h28 == state ? _GEN_96 : iter_ofm_pre; // @[control.scala 438:19 194:31]
  wire [5:0] _GEN_432 = 6'h28 == state ? 6'h29 : _GEN_409; // @[control.scala 1073:19 438:19]
  wire  _GEN_433 = 6'h28 == state ? ifm_send_task_enable : _GEN_408; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_434 = 6'h28 == state ? ifm_addr_fmbase : _GEN_410; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_435 = 6'h28 == state ? ifm_addr_offset : _GEN_411; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_436 = 6'h28 == state ? ifm_send_len : _GEN_412; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_437 = 6'h28 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_413; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_438 = 6'h28 == state ? reg_static : _GEN_414; // @[control.scala 438:19 161:29]
  wire  _GEN_439 = 6'h28 == state ? last_buf_sel : _GEN_415; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_440 = 6'h28 == state ? reg_task : _GEN_416; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_441 = 6'h28 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_417; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_442 = 6'h28 == state ? weight_sel : _GEN_418; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_443 = 6'h28 == state ? wgt_addr_read : _GEN_419; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_444 = 6'h28 == state ? bia_addr_read : _GEN_420; // @[control.scala 438:19 181:32]
  wire  _GEN_445 = 6'h28 == state ? wgt_ddr_read_en : _GEN_421; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_446 = 6'h28 == state ? reg_t_4 : _GEN_422; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_447 = 6'h28 == state ? reg_t_5 : _GEN_423; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_448 = 6'h28 == state ? reg_t_0 : _GEN_424; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_449 = 6'h28 == state ? cnt_t : _GEN_425; // @[control.scala 438:19 163:24]
  wire  _GEN_450 = 6'h28 == state ? ifm_sel : _GEN_426; // @[control.scala 438:19 379:24]
  wire  _GEN_451 = 6'h28 == state ? resize_load_t : _GEN_427; // @[control.scala 438:19 420:32]
  wire  _GEN_452 = 6'h28 == state ? yolo_finish : _GEN_428; // @[control.scala 438:19 40:28]
  wire  _GEN_453 = 6'h28 == state ? conv_finish : _GEN_429; // @[control.scala 438:19 71:30]
  wire  _GEN_454 = 6'h27 == state ? _bottleneck_transfer_T_1 : bottleneck_transfer; // @[control.scala 438:19 1059:33 295:38]
  wire [12:0] _GEN_455 = 6'h27 == state ? _GEN_92 : iter_ifm_pre; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_456 = 6'h27 == state ? _GEN_93 : _GEN_430; // @[control.scala 438:19]
  wire [5:0] _GEN_457 = 6'h27 == state ? _GEN_172 : _GEN_432; // @[control.scala 438:19]
  wire [12:0] _GEN_458 = 6'h27 == state ? iter_ofm_pre : _GEN_431; // @[control.scala 438:19 194:31]
  wire  _GEN_459 = 6'h27 == state ? ifm_send_task_enable : _GEN_433; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_460 = 6'h27 == state ? ifm_addr_fmbase : _GEN_434; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_461 = 6'h27 == state ? ifm_addr_offset : _GEN_435; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_462 = 6'h27 == state ? ifm_send_len : _GEN_436; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_463 = 6'h27 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_437; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_464 = 6'h27 == state ? reg_static : _GEN_438; // @[control.scala 438:19 161:29]
  wire  _GEN_465 = 6'h27 == state ? last_buf_sel : _GEN_439; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_466 = 6'h27 == state ? reg_task : _GEN_440; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_467 = 6'h27 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_441; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_468 = 6'h27 == state ? weight_sel : _GEN_442; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_469 = 6'h27 == state ? wgt_addr_read : _GEN_443; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_470 = 6'h27 == state ? bia_addr_read : _GEN_444; // @[control.scala 438:19 181:32]
  wire  _GEN_471 = 6'h27 == state ? wgt_ddr_read_en : _GEN_445; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_472 = 6'h27 == state ? reg_t_4 : _GEN_446; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_473 = 6'h27 == state ? reg_t_5 : _GEN_447; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_474 = 6'h27 == state ? reg_t_0 : _GEN_448; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_475 = 6'h27 == state ? cnt_t : _GEN_449; // @[control.scala 438:19 163:24]
  wire  _GEN_476 = 6'h27 == state ? ifm_sel : _GEN_450; // @[control.scala 438:19 379:24]
  wire  _GEN_477 = 6'h27 == state ? resize_load_t : _GEN_451; // @[control.scala 438:19 420:32]
  wire  _GEN_478 = 6'h27 == state ? yolo_finish : _GEN_452; // @[control.scala 438:19 40:28]
  wire  _GEN_479 = 6'h27 == state ? conv_finish : _GEN_453; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_480 = 6'h26 == state ? _GEN_165 : _GEN_457; // @[control.scala 438:19]
  wire [12:0] _GEN_481 = 6'h26 == state ? _GEN_166 : iter_ifm_post; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_482 = 6'h26 == state ? _GEN_167 : iter_div_post; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_483 = 6'h26 == state ? _GEN_168 : iter_ofm_post; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_484 = 6'h26 == state ? _GEN_169 : _GEN_455; // @[control.scala 438:19]
  wire  _GEN_485 = 6'h26 == state ? bottleneck_transfer : _GEN_454; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_486 = 6'h26 == state ? iter_div_pre : _GEN_456; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_487 = 6'h26 == state ? iter_ofm_pre : _GEN_458; // @[control.scala 438:19 194:31]
  wire  _GEN_488 = 6'h26 == state ? ifm_send_task_enable : _GEN_459; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_489 = 6'h26 == state ? ifm_addr_fmbase : _GEN_460; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_490 = 6'h26 == state ? ifm_addr_offset : _GEN_461; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_491 = 6'h26 == state ? ifm_send_len : _GEN_462; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_492 = 6'h26 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_463; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_493 = 6'h26 == state ? reg_static : _GEN_464; // @[control.scala 438:19 161:29]
  wire  _GEN_494 = 6'h26 == state ? last_buf_sel : _GEN_465; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_495 = 6'h26 == state ? reg_task : _GEN_466; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_496 = 6'h26 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_467; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_497 = 6'h26 == state ? weight_sel : _GEN_468; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_498 = 6'h26 == state ? wgt_addr_read : _GEN_469; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_499 = 6'h26 == state ? bia_addr_read : _GEN_470; // @[control.scala 438:19 181:32]
  wire  _GEN_500 = 6'h26 == state ? wgt_ddr_read_en : _GEN_471; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_501 = 6'h26 == state ? reg_t_4 : _GEN_472; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_502 = 6'h26 == state ? reg_t_5 : _GEN_473; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_503 = 6'h26 == state ? reg_t_0 : _GEN_474; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_504 = 6'h26 == state ? cnt_t : _GEN_475; // @[control.scala 438:19 163:24]
  wire  _GEN_505 = 6'h26 == state ? ifm_sel : _GEN_476; // @[control.scala 438:19 379:24]
  wire  _GEN_506 = 6'h26 == state ? resize_load_t : _GEN_477; // @[control.scala 438:19 420:32]
  wire  _GEN_507 = 6'h26 == state ? yolo_finish : _GEN_478; // @[control.scala 438:19 40:28]
  wire  _GEN_508 = 6'h26 == state ? conv_finish : _GEN_479; // @[control.scala 438:19 71:30]
  wire [1:0] _GEN_509 = 6'h25 == state ? _GEN_161 : pool_cnt; // @[control.scala 438:19 290:27]
  wire [5:0] _GEN_510 = 6'h25 == state ? _GEN_162 : _GEN_480; // @[control.scala 438:19]
  wire [12:0] _GEN_511 = 6'h25 == state ? iter_ifm_post : _GEN_481; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_512 = 6'h25 == state ? iter_div_post : _GEN_482; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_513 = 6'h25 == state ? iter_ofm_post : _GEN_483; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_514 = 6'h25 == state ? iter_ifm_pre : _GEN_484; // @[control.scala 438:19 192:31]
  wire  _GEN_515 = 6'h25 == state ? bottleneck_transfer : _GEN_485; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_516 = 6'h25 == state ? iter_div_pre : _GEN_486; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_517 = 6'h25 == state ? iter_ofm_pre : _GEN_487; // @[control.scala 438:19 194:31]
  wire  _GEN_518 = 6'h25 == state ? ifm_send_task_enable : _GEN_488; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_519 = 6'h25 == state ? ifm_addr_fmbase : _GEN_489; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_520 = 6'h25 == state ? ifm_addr_offset : _GEN_490; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_521 = 6'h25 == state ? ifm_send_len : _GEN_491; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_522 = 6'h25 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_492; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_523 = 6'h25 == state ? reg_static : _GEN_493; // @[control.scala 438:19 161:29]
  wire  _GEN_524 = 6'h25 == state ? last_buf_sel : _GEN_494; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_525 = 6'h25 == state ? reg_task : _GEN_495; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_526 = 6'h25 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_496; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_527 = 6'h25 == state ? weight_sel : _GEN_497; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_528 = 6'h25 == state ? wgt_addr_read : _GEN_498; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_529 = 6'h25 == state ? bia_addr_read : _GEN_499; // @[control.scala 438:19 181:32]
  wire  _GEN_530 = 6'h25 == state ? wgt_ddr_read_en : _GEN_500; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_531 = 6'h25 == state ? reg_t_4 : _GEN_501; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_532 = 6'h25 == state ? reg_t_5 : _GEN_502; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_533 = 6'h25 == state ? reg_t_0 : _GEN_503; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_534 = 6'h25 == state ? cnt_t : _GEN_504; // @[control.scala 438:19 163:24]
  wire  _GEN_535 = 6'h25 == state ? ifm_sel : _GEN_505; // @[control.scala 438:19 379:24]
  wire  _GEN_536 = 6'h25 == state ? resize_load_t : _GEN_506; // @[control.scala 438:19 420:32]
  wire  _GEN_537 = 6'h25 == state ? yolo_finish : _GEN_507; // @[control.scala 438:19 40:28]
  wire  _GEN_538 = 6'h25 == state ? conv_finish : _GEN_508; // @[control.scala 438:19 71:30]
  wire [4:0] _GEN_539 = 6'h24 == state ? _GEN_2 : _GEN_534; // @[control.scala 438:19]
  wire [31:0] _GEN_540 = 6'h24 == state ? _GEN_71 : _GEN_533; // @[control.scala 438:19]
  wire [5:0] _GEN_541 = 6'h24 == state ? _GEN_156 : _GEN_510; // @[control.scala 438:19]
  wire [1:0] _GEN_542 = 6'h24 == state ? pool_cnt : _GEN_509; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_543 = 6'h24 == state ? iter_ifm_post : _GEN_511; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_544 = 6'h24 == state ? iter_div_post : _GEN_512; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_545 = 6'h24 == state ? iter_ofm_post : _GEN_513; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_546 = 6'h24 == state ? iter_ifm_pre : _GEN_514; // @[control.scala 438:19 192:31]
  wire  _GEN_547 = 6'h24 == state ? bottleneck_transfer : _GEN_515; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_548 = 6'h24 == state ? iter_div_pre : _GEN_516; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_549 = 6'h24 == state ? iter_ofm_pre : _GEN_517; // @[control.scala 438:19 194:31]
  wire  _GEN_550 = 6'h24 == state ? ifm_send_task_enable : _GEN_518; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_551 = 6'h24 == state ? ifm_addr_fmbase : _GEN_519; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_552 = 6'h24 == state ? ifm_addr_offset : _GEN_520; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_553 = 6'h24 == state ? ifm_send_len : _GEN_521; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_554 = 6'h24 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_522; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_555 = 6'h24 == state ? reg_static : _GEN_523; // @[control.scala 438:19 161:29]
  wire  _GEN_556 = 6'h24 == state ? last_buf_sel : _GEN_524; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_557 = 6'h24 == state ? reg_task : _GEN_525; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_558 = 6'h24 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_526; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_559 = 6'h24 == state ? weight_sel : _GEN_527; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_560 = 6'h24 == state ? wgt_addr_read : _GEN_528; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_561 = 6'h24 == state ? bia_addr_read : _GEN_529; // @[control.scala 438:19 181:32]
  wire  _GEN_562 = 6'h24 == state ? wgt_ddr_read_en : _GEN_530; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_563 = 6'h24 == state ? reg_t_4 : _GEN_531; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_564 = 6'h24 == state ? reg_t_5 : _GEN_532; // @[control.scala 438:19 160:37]
  wire  _GEN_565 = 6'h24 == state ? ifm_sel : _GEN_535; // @[control.scala 438:19 379:24]
  wire  _GEN_566 = 6'h24 == state ? resize_load_t : _GEN_536; // @[control.scala 438:19 420:32]
  wire  _GEN_567 = 6'h24 == state ? yolo_finish : _GEN_537; // @[control.scala 438:19 40:28]
  wire  _GEN_568 = 6'h24 == state ? conv_finish : _GEN_538; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_569 = 6'h23 == state ? ofm_addr_recv : reg_t_6; // @[control.scala 438:19 1002:22 160:37]
  wire [31:0] _GEN_570 = 6'h23 == state ? ofm_recv_len : reg_t_7; // @[control.scala 438:19 1003:22 160:37]
  wire [31:0] _GEN_571 = 6'h23 == state ? _reg_t_0_T_7 : _GEN_540; // @[control.scala 438:19 1005:22]
  wire [4:0] _GEN_572 = 6'h23 == state ? 5'h0 : _GEN_539; // @[control.scala 1006:19 438:19]
  wire [5:0] _GEN_573 = 6'h23 == state ? 6'h24 : _GEN_541; // @[control.scala 1007:19 438:19]
  wire [1:0] _GEN_574 = 6'h23 == state ? pool_cnt : _GEN_542; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_575 = 6'h23 == state ? iter_ifm_post : _GEN_543; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_576 = 6'h23 == state ? iter_div_post : _GEN_544; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_577 = 6'h23 == state ? iter_ofm_post : _GEN_545; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_578 = 6'h23 == state ? iter_ifm_pre : _GEN_546; // @[control.scala 438:19 192:31]
  wire  _GEN_579 = 6'h23 == state ? bottleneck_transfer : _GEN_547; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_580 = 6'h23 == state ? iter_div_pre : _GEN_548; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_581 = 6'h23 == state ? iter_ofm_pre : _GEN_549; // @[control.scala 438:19 194:31]
  wire  _GEN_582 = 6'h23 == state ? ifm_send_task_enable : _GEN_550; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_583 = 6'h23 == state ? ifm_addr_fmbase : _GEN_551; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_584 = 6'h23 == state ? ifm_addr_offset : _GEN_552; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_585 = 6'h23 == state ? ifm_send_len : _GEN_553; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_586 = 6'h23 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_554; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_587 = 6'h23 == state ? reg_static : _GEN_555; // @[control.scala 438:19 161:29]
  wire  _GEN_588 = 6'h23 == state ? last_buf_sel : _GEN_556; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_589 = 6'h23 == state ? reg_task : _GEN_557; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_590 = 6'h23 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_558; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_591 = 6'h23 == state ? weight_sel : _GEN_559; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_592 = 6'h23 == state ? wgt_addr_read : _GEN_560; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_593 = 6'h23 == state ? bia_addr_read : _GEN_561; // @[control.scala 438:19 181:32]
  wire  _GEN_594 = 6'h23 == state ? wgt_ddr_read_en : _GEN_562; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_595 = 6'h23 == state ? reg_t_4 : _GEN_563; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_596 = 6'h23 == state ? reg_t_5 : _GEN_564; // @[control.scala 438:19 160:37]
  wire  _GEN_597 = 6'h23 == state ? ifm_sel : _GEN_565; // @[control.scala 438:19 379:24]
  wire  _GEN_598 = 6'h23 == state ? resize_load_t : _GEN_566; // @[control.scala 438:19 420:32]
  wire  _GEN_599 = 6'h23 == state ? yolo_finish : _GEN_567; // @[control.scala 438:19 40:28]
  wire  _GEN_600 = 6'h23 == state ? conv_finish : _GEN_568; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_601 = 6'h22 == state ? _GEN_154 : _GEN_573; // @[control.scala 438:19]
  wire [31:0] _GEN_602 = 6'h22 == state ? reg_t_6 : _GEN_569; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_603 = 6'h22 == state ? reg_t_7 : _GEN_570; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_604 = 6'h22 == state ? reg_t_0 : _GEN_571; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_605 = 6'h22 == state ? cnt_t : _GEN_572; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_606 = 6'h22 == state ? pool_cnt : _GEN_574; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_607 = 6'h22 == state ? iter_ifm_post : _GEN_575; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_608 = 6'h22 == state ? iter_div_post : _GEN_576; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_609 = 6'h22 == state ? iter_ofm_post : _GEN_577; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_610 = 6'h22 == state ? iter_ifm_pre : _GEN_578; // @[control.scala 438:19 192:31]
  wire  _GEN_611 = 6'h22 == state ? bottleneck_transfer : _GEN_579; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_612 = 6'h22 == state ? iter_div_pre : _GEN_580; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_613 = 6'h22 == state ? iter_ofm_pre : _GEN_581; // @[control.scala 438:19 194:31]
  wire  _GEN_614 = 6'h22 == state ? ifm_send_task_enable : _GEN_582; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_615 = 6'h22 == state ? ifm_addr_fmbase : _GEN_583; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_616 = 6'h22 == state ? ifm_addr_offset : _GEN_584; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_617 = 6'h22 == state ? ifm_send_len : _GEN_585; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_618 = 6'h22 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_586; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_619 = 6'h22 == state ? reg_static : _GEN_587; // @[control.scala 438:19 161:29]
  wire  _GEN_620 = 6'h22 == state ? last_buf_sel : _GEN_588; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_621 = 6'h22 == state ? reg_task : _GEN_589; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_622 = 6'h22 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_590; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_623 = 6'h22 == state ? weight_sel : _GEN_591; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_624 = 6'h22 == state ? wgt_addr_read : _GEN_592; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_625 = 6'h22 == state ? bia_addr_read : _GEN_593; // @[control.scala 438:19 181:32]
  wire  _GEN_626 = 6'h22 == state ? wgt_ddr_read_en : _GEN_594; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_627 = 6'h22 == state ? reg_t_4 : _GEN_595; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_628 = 6'h22 == state ? reg_t_5 : _GEN_596; // @[control.scala 438:19 160:37]
  wire  _GEN_629 = 6'h22 == state ? ifm_sel : _GEN_597; // @[control.scala 438:19 379:24]
  wire  _GEN_630 = 6'h22 == state ? resize_load_t : _GEN_598; // @[control.scala 438:19 420:32]
  wire  _GEN_631 = 6'h22 == state ? yolo_finish : _GEN_599; // @[control.scala 438:19 40:28]
  wire  _GEN_632 = 6'h22 == state ? conv_finish : _GEN_600; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_633 = 6'h21 == state ? _reg_t_0_T_5 : _GEN_604; // @[control.scala 438:19 987:22]
  wire [5:0] _GEN_634 = 6'h21 == state ? 6'h22 : _GEN_601; // @[control.scala 438:19 988:19]
  wire [31:0] _GEN_635 = 6'h21 == state ? reg_t_6 : _GEN_602; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_636 = 6'h21 == state ? reg_t_7 : _GEN_603; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_637 = 6'h21 == state ? cnt_t : _GEN_605; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_638 = 6'h21 == state ? pool_cnt : _GEN_606; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_639 = 6'h21 == state ? iter_ifm_post : _GEN_607; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_640 = 6'h21 == state ? iter_div_post : _GEN_608; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_641 = 6'h21 == state ? iter_ofm_post : _GEN_609; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_642 = 6'h21 == state ? iter_ifm_pre : _GEN_610; // @[control.scala 438:19 192:31]
  wire  _GEN_643 = 6'h21 == state ? bottleneck_transfer : _GEN_611; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_644 = 6'h21 == state ? iter_div_pre : _GEN_612; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_645 = 6'h21 == state ? iter_ofm_pre : _GEN_613; // @[control.scala 438:19 194:31]
  wire  _GEN_646 = 6'h21 == state ? ifm_send_task_enable : _GEN_614; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_647 = 6'h21 == state ? ifm_addr_fmbase : _GEN_615; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_648 = 6'h21 == state ? ifm_addr_offset : _GEN_616; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_649 = 6'h21 == state ? ifm_send_len : _GEN_617; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_650 = 6'h21 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_618; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_651 = 6'h21 == state ? reg_static : _GEN_619; // @[control.scala 438:19 161:29]
  wire  _GEN_652 = 6'h21 == state ? last_buf_sel : _GEN_620; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_653 = 6'h21 == state ? reg_task : _GEN_621; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_654 = 6'h21 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_622; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_655 = 6'h21 == state ? weight_sel : _GEN_623; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_656 = 6'h21 == state ? wgt_addr_read : _GEN_624; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_657 = 6'h21 == state ? bia_addr_read : _GEN_625; // @[control.scala 438:19 181:32]
  wire  _GEN_658 = 6'h21 == state ? wgt_ddr_read_en : _GEN_626; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_659 = 6'h21 == state ? reg_t_4 : _GEN_627; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_660 = 6'h21 == state ? reg_t_5 : _GEN_628; // @[control.scala 438:19 160:37]
  wire  _GEN_661 = 6'h21 == state ? ifm_sel : _GEN_629; // @[control.scala 438:19 379:24]
  wire  _GEN_662 = 6'h21 == state ? resize_load_t : _GEN_630; // @[control.scala 438:19 420:32]
  wire  _GEN_663 = 6'h21 == state ? yolo_finish : _GEN_631; // @[control.scala 438:19 40:28]
  wire  _GEN_664 = 6'h21 == state ? conv_finish : _GEN_632; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_665 = 6'h20 == state ? _GEN_153 : _GEN_634; // @[control.scala 438:19]
  wire [31:0] _GEN_666 = 6'h20 == state ? reg_t_0 : _GEN_633; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_667 = 6'h20 == state ? reg_t_6 : _GEN_635; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_668 = 6'h20 == state ? reg_t_7 : _GEN_636; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_669 = 6'h20 == state ? cnt_t : _GEN_637; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_670 = 6'h20 == state ? pool_cnt : _GEN_638; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_671 = 6'h20 == state ? iter_ifm_post : _GEN_639; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_672 = 6'h20 == state ? iter_div_post : _GEN_640; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_673 = 6'h20 == state ? iter_ofm_post : _GEN_641; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_674 = 6'h20 == state ? iter_ifm_pre : _GEN_642; // @[control.scala 438:19 192:31]
  wire  _GEN_675 = 6'h20 == state ? bottleneck_transfer : _GEN_643; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_676 = 6'h20 == state ? iter_div_pre : _GEN_644; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_677 = 6'h20 == state ? iter_ofm_pre : _GEN_645; // @[control.scala 438:19 194:31]
  wire  _GEN_678 = 6'h20 == state ? ifm_send_task_enable : _GEN_646; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_679 = 6'h20 == state ? ifm_addr_fmbase : _GEN_647; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_680 = 6'h20 == state ? ifm_addr_offset : _GEN_648; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_681 = 6'h20 == state ? ifm_send_len : _GEN_649; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_682 = 6'h20 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_650; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_683 = 6'h20 == state ? reg_static : _GEN_651; // @[control.scala 438:19 161:29]
  wire  _GEN_684 = 6'h20 == state ? last_buf_sel : _GEN_652; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_685 = 6'h20 == state ? reg_task : _GEN_653; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_686 = 6'h20 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_654; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_687 = 6'h20 == state ? weight_sel : _GEN_655; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_688 = 6'h20 == state ? wgt_addr_read : _GEN_656; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_689 = 6'h20 == state ? bia_addr_read : _GEN_657; // @[control.scala 438:19 181:32]
  wire  _GEN_690 = 6'h20 == state ? wgt_ddr_read_en : _GEN_658; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_691 = 6'h20 == state ? reg_t_4 : _GEN_659; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_692 = 6'h20 == state ? reg_t_5 : _GEN_660; // @[control.scala 438:19 160:37]
  wire  _GEN_693 = 6'h20 == state ? ifm_sel : _GEN_661; // @[control.scala 438:19 379:24]
  wire  _GEN_694 = 6'h20 == state ? resize_load_t : _GEN_662; // @[control.scala 438:19 420:32]
  wire  _GEN_695 = 6'h20 == state ? yolo_finish : _GEN_663; // @[control.scala 438:19 40:28]
  wire  _GEN_696 = 6'h20 == state ? conv_finish : _GEN_664; // @[control.scala 438:19 71:30]
  wire [15:0] _GEN_697 = 6'h1f == state ? _wgt_addr_read_T : _GEN_688; // @[control.scala 438:19 967:27]
  wire [15:0] _GEN_698 = 6'h1f == state ? {{3'd0}, iter_ofm_post} : _GEN_689; // @[control.scala 438:19 968:27]
  wire  _GEN_699 = 6'h1f == state ? _wgt_ddr_read_en_T_6 : _GEN_690; // @[control.scala 438:19 969:28]
  wire [5:0] _GEN_700 = 6'h1f == state ? 6'h20 : _GEN_665; // @[control.scala 438:19 970:19]
  wire [31:0] _GEN_701 = 6'h1f == state ? reg_t_0 : _GEN_666; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_702 = 6'h1f == state ? reg_t_6 : _GEN_667; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_703 = 6'h1f == state ? reg_t_7 : _GEN_668; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_704 = 6'h1f == state ? cnt_t : _GEN_669; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_705 = 6'h1f == state ? pool_cnt : _GEN_670; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_706 = 6'h1f == state ? iter_ifm_post : _GEN_671; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_707 = 6'h1f == state ? iter_div_post : _GEN_672; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_708 = 6'h1f == state ? iter_ofm_post : _GEN_673; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_709 = 6'h1f == state ? iter_ifm_pre : _GEN_674; // @[control.scala 438:19 192:31]
  wire  _GEN_710 = 6'h1f == state ? bottleneck_transfer : _GEN_675; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_711 = 6'h1f == state ? iter_div_pre : _GEN_676; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_712 = 6'h1f == state ? iter_ofm_pre : _GEN_677; // @[control.scala 438:19 194:31]
  wire  _GEN_713 = 6'h1f == state ? ifm_send_task_enable : _GEN_678; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_714 = 6'h1f == state ? ifm_addr_fmbase : _GEN_679; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_715 = 6'h1f == state ? ifm_addr_offset : _GEN_680; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_716 = 6'h1f == state ? ifm_send_len : _GEN_681; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_717 = 6'h1f == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_682; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_718 = 6'h1f == state ? reg_static : _GEN_683; // @[control.scala 438:19 161:29]
  wire  _GEN_719 = 6'h1f == state ? last_buf_sel : _GEN_684; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_720 = 6'h1f == state ? reg_task : _GEN_685; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_721 = 6'h1f == state ? {{10'd0}, wgt_addr_read_t} : _GEN_686; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_722 = 6'h1f == state ? weight_sel : _GEN_687; // @[control.scala 438:19 274:27]
  wire [31:0] _GEN_723 = 6'h1f == state ? reg_t_4 : _GEN_691; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_724 = 6'h1f == state ? reg_t_5 : _GEN_692; // @[control.scala 438:19 160:37]
  wire  _GEN_725 = 6'h1f == state ? ifm_sel : _GEN_693; // @[control.scala 438:19 379:24]
  wire  _GEN_726 = 6'h1f == state ? resize_load_t : _GEN_694; // @[control.scala 438:19 420:32]
  wire  _GEN_727 = 6'h1f == state ? yolo_finish : _GEN_695; // @[control.scala 438:19 40:28]
  wire  _GEN_728 = 6'h1f == state ? conv_finish : _GEN_696; // @[control.scala 438:19 71:30]
  wire [25:0] _GEN_729 = 6'h1e == state ? _GEN_150 : _GEN_721; // @[control.scala 438:19]
  wire [2:0] _GEN_730 = 6'h1e == state ? _GEN_151 : _GEN_722; // @[control.scala 438:19]
  wire [5:0] _GEN_731 = 6'h1e == state ? 6'h1f : _GEN_700; // @[control.scala 438:19 964:19]
  wire [15:0] _GEN_732 = 6'h1e == state ? wgt_addr_read : _GEN_697; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_733 = 6'h1e == state ? bia_addr_read : _GEN_698; // @[control.scala 438:19 181:32]
  wire  _GEN_734 = 6'h1e == state ? wgt_ddr_read_en : _GEN_699; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_735 = 6'h1e == state ? reg_t_0 : _GEN_701; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_736 = 6'h1e == state ? reg_t_6 : _GEN_702; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_737 = 6'h1e == state ? reg_t_7 : _GEN_703; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_738 = 6'h1e == state ? cnt_t : _GEN_704; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_739 = 6'h1e == state ? pool_cnt : _GEN_705; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_740 = 6'h1e == state ? iter_ifm_post : _GEN_706; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_741 = 6'h1e == state ? iter_div_post : _GEN_707; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_742 = 6'h1e == state ? iter_ofm_post : _GEN_708; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_743 = 6'h1e == state ? iter_ifm_pre : _GEN_709; // @[control.scala 438:19 192:31]
  wire  _GEN_744 = 6'h1e == state ? bottleneck_transfer : _GEN_710; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_745 = 6'h1e == state ? iter_div_pre : _GEN_711; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_746 = 6'h1e == state ? iter_ofm_pre : _GEN_712; // @[control.scala 438:19 194:31]
  wire  _GEN_747 = 6'h1e == state ? ifm_send_task_enable : _GEN_713; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_748 = 6'h1e == state ? ifm_addr_fmbase : _GEN_714; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_749 = 6'h1e == state ? ifm_addr_offset : _GEN_715; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_750 = 6'h1e == state ? ifm_send_len : _GEN_716; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_751 = 6'h1e == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_717; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_752 = 6'h1e == state ? reg_static : _GEN_718; // @[control.scala 438:19 161:29]
  wire  _GEN_753 = 6'h1e == state ? last_buf_sel : _GEN_719; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_754 = 6'h1e == state ? reg_task : _GEN_720; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_755 = 6'h1e == state ? reg_t_4 : _GEN_723; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_756 = 6'h1e == state ? reg_t_5 : _GEN_724; // @[control.scala 438:19 160:37]
  wire  _GEN_757 = 6'h1e == state ? ifm_sel : _GEN_725; // @[control.scala 438:19 379:24]
  wire  _GEN_758 = 6'h1e == state ? resize_load_t : _GEN_726; // @[control.scala 438:19 420:32]
  wire  _GEN_759 = 6'h1e == state ? yolo_finish : _GEN_727; // @[control.scala 438:19 40:28]
  wire  _GEN_760 = 6'h1e == state ? conv_finish : _GEN_728; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_761 = 6'h1d == state ? _GEN_62 : _GEN_752; // @[control.scala 438:19]
  wire [31:0] _GEN_762 = 6'h1d == state ? {{22'd0}, _GEN_148} : _GEN_754; // @[control.scala 438:19]
  wire [5:0] _GEN_763 = 6'h1d == state ? 6'h1e : _GEN_731; // @[control.scala 438:19 950:19]
  wire [25:0] _GEN_764 = 6'h1d == state ? {{10'd0}, wgt_addr_read_t} : _GEN_729; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_765 = 6'h1d == state ? weight_sel : _GEN_730; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_766 = 6'h1d == state ? wgt_addr_read : _GEN_732; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_767 = 6'h1d == state ? bia_addr_read : _GEN_733; // @[control.scala 438:19 181:32]
  wire  _GEN_768 = 6'h1d == state ? wgt_ddr_read_en : _GEN_734; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_769 = 6'h1d == state ? reg_t_0 : _GEN_735; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_770 = 6'h1d == state ? reg_t_6 : _GEN_736; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_771 = 6'h1d == state ? reg_t_7 : _GEN_737; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_772 = 6'h1d == state ? cnt_t : _GEN_738; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_773 = 6'h1d == state ? pool_cnt : _GEN_739; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_774 = 6'h1d == state ? iter_ifm_post : _GEN_740; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_775 = 6'h1d == state ? iter_div_post : _GEN_741; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_776 = 6'h1d == state ? iter_ofm_post : _GEN_742; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_777 = 6'h1d == state ? iter_ifm_pre : _GEN_743; // @[control.scala 438:19 192:31]
  wire  _GEN_778 = 6'h1d == state ? bottleneck_transfer : _GEN_744; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_779 = 6'h1d == state ? iter_div_pre : _GEN_745; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_780 = 6'h1d == state ? iter_ofm_pre : _GEN_746; // @[control.scala 438:19 194:31]
  wire  _GEN_781 = 6'h1d == state ? ifm_send_task_enable : _GEN_747; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_782 = 6'h1d == state ? ifm_addr_fmbase : _GEN_748; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_783 = 6'h1d == state ? ifm_addr_offset : _GEN_749; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_784 = 6'h1d == state ? ifm_send_len : _GEN_750; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_785 = 6'h1d == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_751; // @[control.scala 438:19 425:46]
  wire  _GEN_786 = 6'h1d == state ? last_buf_sel : _GEN_753; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_787 = 6'h1d == state ? reg_t_4 : _GEN_755; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_788 = 6'h1d == state ? reg_t_5 : _GEN_756; // @[control.scala 438:19 160:37]
  wire  _GEN_789 = 6'h1d == state ? ifm_sel : _GEN_757; // @[control.scala 438:19 379:24]
  wire  _GEN_790 = 6'h1d == state ? resize_load_t : _GEN_758; // @[control.scala 438:19 420:32]
  wire  _GEN_791 = 6'h1d == state ? yolo_finish : _GEN_759; // @[control.scala 438:19 40:28]
  wire  _GEN_792 = 6'h1d == state ? conv_finish : _GEN_760; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_793 = 6'h1c == state ? _GEN_55 : _GEN_761; // @[control.scala 438:19]
  wire [5:0] _GEN_794 = 6'h1c == state ? 6'h1d : _GEN_763; // @[control.scala 438:19 912:18]
  wire [31:0] _GEN_795 = 6'h1c == state ? reg_task : _GEN_762; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_796 = 6'h1c == state ? {{10'd0}, wgt_addr_read_t} : _GEN_764; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_797 = 6'h1c == state ? weight_sel : _GEN_765; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_798 = 6'h1c == state ? wgt_addr_read : _GEN_766; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_799 = 6'h1c == state ? bia_addr_read : _GEN_767; // @[control.scala 438:19 181:32]
  wire  _GEN_800 = 6'h1c == state ? wgt_ddr_read_en : _GEN_768; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_801 = 6'h1c == state ? reg_t_0 : _GEN_769; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_802 = 6'h1c == state ? reg_t_6 : _GEN_770; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_803 = 6'h1c == state ? reg_t_7 : _GEN_771; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_804 = 6'h1c == state ? cnt_t : _GEN_772; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_805 = 6'h1c == state ? pool_cnt : _GEN_773; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_806 = 6'h1c == state ? iter_ifm_post : _GEN_774; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_807 = 6'h1c == state ? iter_div_post : _GEN_775; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_808 = 6'h1c == state ? iter_ofm_post : _GEN_776; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_809 = 6'h1c == state ? iter_ifm_pre : _GEN_777; // @[control.scala 438:19 192:31]
  wire  _GEN_810 = 6'h1c == state ? bottleneck_transfer : _GEN_778; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_811 = 6'h1c == state ? iter_div_pre : _GEN_779; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_812 = 6'h1c == state ? iter_ofm_pre : _GEN_780; // @[control.scala 438:19 194:31]
  wire  _GEN_813 = 6'h1c == state ? ifm_send_task_enable : _GEN_781; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_814 = 6'h1c == state ? ifm_addr_fmbase : _GEN_782; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_815 = 6'h1c == state ? ifm_addr_offset : _GEN_783; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_816 = 6'h1c == state ? ifm_send_len : _GEN_784; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_817 = 6'h1c == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_785; // @[control.scala 438:19 425:46]
  wire  _GEN_818 = 6'h1c == state ? last_buf_sel : _GEN_786; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_819 = 6'h1c == state ? reg_t_4 : _GEN_787; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_820 = 6'h1c == state ? reg_t_5 : _GEN_788; // @[control.scala 438:19 160:37]
  wire  _GEN_821 = 6'h1c == state ? ifm_sel : _GEN_789; // @[control.scala 438:19 379:24]
  wire  _GEN_822 = 6'h1c == state ? resize_load_t : _GEN_790; // @[control.scala 438:19 420:32]
  wire  _GEN_823 = 6'h1c == state ? yolo_finish : _GEN_791; // @[control.scala 438:19 40:28]
  wire  _GEN_824 = 6'h1c == state ? conv_finish : _GEN_792; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_825 = 6'h1b == state ? _GEN_52 : _GEN_793; // @[control.scala 438:19]
  wire  _GEN_826 = 6'h1b == state ? _T_28 : _GEN_818; // @[control.scala 438:19 901:26]
  wire [5:0] _GEN_827 = 6'h1b == state ? 6'h1c : _GEN_794; // @[control.scala 438:19 902:19]
  wire [31:0] _GEN_828 = 6'h1b == state ? reg_task : _GEN_795; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_829 = 6'h1b == state ? {{10'd0}, wgt_addr_read_t} : _GEN_796; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_830 = 6'h1b == state ? weight_sel : _GEN_797; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_831 = 6'h1b == state ? wgt_addr_read : _GEN_798; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_832 = 6'h1b == state ? bia_addr_read : _GEN_799; // @[control.scala 438:19 181:32]
  wire  _GEN_833 = 6'h1b == state ? wgt_ddr_read_en : _GEN_800; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_834 = 6'h1b == state ? reg_t_0 : _GEN_801; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_835 = 6'h1b == state ? reg_t_6 : _GEN_802; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_836 = 6'h1b == state ? reg_t_7 : _GEN_803; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_837 = 6'h1b == state ? cnt_t : _GEN_804; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_838 = 6'h1b == state ? pool_cnt : _GEN_805; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_839 = 6'h1b == state ? iter_ifm_post : _GEN_806; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_840 = 6'h1b == state ? iter_div_post : _GEN_807; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_841 = 6'h1b == state ? iter_ofm_post : _GEN_808; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_842 = 6'h1b == state ? iter_ifm_pre : _GEN_809; // @[control.scala 438:19 192:31]
  wire  _GEN_843 = 6'h1b == state ? bottleneck_transfer : _GEN_810; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_844 = 6'h1b == state ? iter_div_pre : _GEN_811; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_845 = 6'h1b == state ? iter_ofm_pre : _GEN_812; // @[control.scala 438:19 194:31]
  wire  _GEN_846 = 6'h1b == state ? ifm_send_task_enable : _GEN_813; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_847 = 6'h1b == state ? ifm_addr_fmbase : _GEN_814; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_848 = 6'h1b == state ? ifm_addr_offset : _GEN_815; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_849 = 6'h1b == state ? ifm_send_len : _GEN_816; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_850 = 6'h1b == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_817; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_851 = 6'h1b == state ? reg_t_4 : _GEN_819; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_852 = 6'h1b == state ? reg_t_5 : _GEN_820; // @[control.scala 438:19 160:37]
  wire  _GEN_853 = 6'h1b == state ? ifm_sel : _GEN_821; // @[control.scala 438:19 379:24]
  wire  _GEN_854 = 6'h1b == state ? resize_load_t : _GEN_822; // @[control.scala 438:19 420:32]
  wire  _GEN_855 = 6'h1b == state ? yolo_finish : _GEN_823; // @[control.scala 438:19 40:28]
  wire  _GEN_856 = 6'h1b == state ? conv_finish : _GEN_824; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_857 = 6'h1a == state ? _GEN_51 : _GEN_825; // @[control.scala 438:19]
  wire [5:0] _GEN_858 = 6'h1a == state ? 6'h1b : _GEN_827; // @[control.scala 438:19 894:19]
  wire  _GEN_859 = 6'h1a == state ? last_buf_sel : _GEN_826; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_860 = 6'h1a == state ? reg_task : _GEN_828; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_861 = 6'h1a == state ? {{10'd0}, wgt_addr_read_t} : _GEN_829; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_862 = 6'h1a == state ? weight_sel : _GEN_830; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_863 = 6'h1a == state ? wgt_addr_read : _GEN_831; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_864 = 6'h1a == state ? bia_addr_read : _GEN_832; // @[control.scala 438:19 181:32]
  wire  _GEN_865 = 6'h1a == state ? wgt_ddr_read_en : _GEN_833; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_866 = 6'h1a == state ? reg_t_0 : _GEN_834; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_867 = 6'h1a == state ? reg_t_6 : _GEN_835; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_868 = 6'h1a == state ? reg_t_7 : _GEN_836; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_869 = 6'h1a == state ? cnt_t : _GEN_837; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_870 = 6'h1a == state ? pool_cnt : _GEN_838; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_871 = 6'h1a == state ? iter_ifm_post : _GEN_839; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_872 = 6'h1a == state ? iter_div_post : _GEN_840; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_873 = 6'h1a == state ? iter_ofm_post : _GEN_841; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_874 = 6'h1a == state ? iter_ifm_pre : _GEN_842; // @[control.scala 438:19 192:31]
  wire  _GEN_875 = 6'h1a == state ? bottleneck_transfer : _GEN_843; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_876 = 6'h1a == state ? iter_div_pre : _GEN_844; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_877 = 6'h1a == state ? iter_ofm_pre : _GEN_845; // @[control.scala 438:19 194:31]
  wire  _GEN_878 = 6'h1a == state ? ifm_send_task_enable : _GEN_846; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_879 = 6'h1a == state ? ifm_addr_fmbase : _GEN_847; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_880 = 6'h1a == state ? ifm_addr_offset : _GEN_848; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_881 = 6'h1a == state ? ifm_send_len : _GEN_849; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_882 = 6'h1a == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_850; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_883 = 6'h1a == state ? reg_t_4 : _GEN_851; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_884 = 6'h1a == state ? reg_t_5 : _GEN_852; // @[control.scala 438:19 160:37]
  wire  _GEN_885 = 6'h1a == state ? ifm_sel : _GEN_853; // @[control.scala 438:19 379:24]
  wire  _GEN_886 = 6'h1a == state ? resize_load_t : _GEN_854; // @[control.scala 438:19 420:32]
  wire  _GEN_887 = 6'h1a == state ? yolo_finish : _GEN_855; // @[control.scala 438:19 40:28]
  wire  _GEN_888 = 6'h1a == state ? conv_finish : _GEN_856; // @[control.scala 438:19 71:30]
  wire  _GEN_889 = 6'h19 == state | _GEN_878; // @[control.scala 438:19 866:34]
  wire [31:0] _GEN_890 = 6'h19 == state ? _ofm_addr_fmbase_T : _GEN_879; // @[control.scala 438:19 867:29]
  wire [31:0] _GEN_891 = 6'h19 == state ? _GEN_131 : _GEN_880; // @[control.scala 438:19]
  wire [31:0] _GEN_892 = 6'h19 == state ? {{10'd0}, _GEN_132} : _GEN_881; // @[control.scala 438:19]
  wire [5:0] _GEN_893 = 6'h19 == state ? 6'h1a : _GEN_858; // @[control.scala 438:19 880:19]
  wire [31:0] _GEN_894 = 6'h19 == state ? reg_static : _GEN_857; // @[control.scala 438:19 161:29]
  wire  _GEN_895 = 6'h19 == state ? last_buf_sel : _GEN_859; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_896 = 6'h19 == state ? reg_task : _GEN_860; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_897 = 6'h19 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_861; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_898 = 6'h19 == state ? weight_sel : _GEN_862; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_899 = 6'h19 == state ? wgt_addr_read : _GEN_863; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_900 = 6'h19 == state ? bia_addr_read : _GEN_864; // @[control.scala 438:19 181:32]
  wire  _GEN_901 = 6'h19 == state ? wgt_ddr_read_en : _GEN_865; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_902 = 6'h19 == state ? reg_t_0 : _GEN_866; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_903 = 6'h19 == state ? reg_t_6 : _GEN_867; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_904 = 6'h19 == state ? reg_t_7 : _GEN_868; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_905 = 6'h19 == state ? cnt_t : _GEN_869; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_906 = 6'h19 == state ? pool_cnt : _GEN_870; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_907 = 6'h19 == state ? iter_ifm_post : _GEN_871; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_908 = 6'h19 == state ? iter_div_post : _GEN_872; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_909 = 6'h19 == state ? iter_ofm_post : _GEN_873; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_910 = 6'h19 == state ? iter_ifm_pre : _GEN_874; // @[control.scala 438:19 192:31]
  wire  _GEN_911 = 6'h19 == state ? bottleneck_transfer : _GEN_875; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_912 = 6'h19 == state ? iter_div_pre : _GEN_876; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_913 = 6'h19 == state ? iter_ofm_pre : _GEN_877; // @[control.scala 438:19 194:31]
  wire [9:0] _GEN_914 = 6'h19 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_882; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_915 = 6'h19 == state ? reg_t_4 : _GEN_883; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_916 = 6'h19 == state ? reg_t_5 : _GEN_884; // @[control.scala 438:19 160:37]
  wire  _GEN_917 = 6'h19 == state ? ifm_sel : _GEN_885; // @[control.scala 438:19 379:24]
  wire  _GEN_918 = 6'h19 == state ? resize_load_t : _GEN_886; // @[control.scala 438:19 420:32]
  wire  _GEN_919 = 6'h19 == state ? yolo_finish : _GEN_887; // @[control.scala 438:19 40:28]
  wire  _GEN_920 = 6'h19 == state ? conv_finish : _GEN_888; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_921 = 6'h18 == state ? _ifm_addr_fmbase_T : _GEN_890; // @[control.scala 438:19 811:29]
  wire [31:0] _GEN_922 = 6'h18 == state ? _GEN_45 : _GEN_891; // @[control.scala 438:19]
  wire [31:0] _GEN_923 = 6'h18 == state ? _GEN_46 : _GEN_892; // @[control.scala 438:19]
  wire [9:0] _GEN_924 = 6'h18 == state ? _GEN_47 : _GEN_914; // @[control.scala 438:19]
  wire [31:0] _GEN_925 = 6'h18 == state ? _GEN_48 : _GEN_894; // @[control.scala 438:19]
  wire [5:0] _GEN_926 = 6'h18 == state ? 6'h1a : _GEN_893; // @[control.scala 438:19 863:19]
  wire  _GEN_927 = 6'h18 == state ? ifm_send_task_enable : _GEN_889; // @[control.scala 438:19 357:39]
  wire  _GEN_928 = 6'h18 == state ? last_buf_sel : _GEN_895; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_929 = 6'h18 == state ? reg_task : _GEN_896; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_930 = 6'h18 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_897; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_931 = 6'h18 == state ? weight_sel : _GEN_898; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_932 = 6'h18 == state ? wgt_addr_read : _GEN_899; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_933 = 6'h18 == state ? bia_addr_read : _GEN_900; // @[control.scala 438:19 181:32]
  wire  _GEN_934 = 6'h18 == state ? wgt_ddr_read_en : _GEN_901; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_935 = 6'h18 == state ? reg_t_0 : _GEN_902; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_936 = 6'h18 == state ? reg_t_6 : _GEN_903; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_937 = 6'h18 == state ? reg_t_7 : _GEN_904; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_938 = 6'h18 == state ? cnt_t : _GEN_905; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_939 = 6'h18 == state ? pool_cnt : _GEN_906; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_940 = 6'h18 == state ? iter_ifm_post : _GEN_907; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_941 = 6'h18 == state ? iter_div_post : _GEN_908; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_942 = 6'h18 == state ? iter_ofm_post : _GEN_909; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_943 = 6'h18 == state ? iter_ifm_pre : _GEN_910; // @[control.scala 438:19 192:31]
  wire  _GEN_944 = 6'h18 == state ? bottleneck_transfer : _GEN_911; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_945 = 6'h18 == state ? iter_div_pre : _GEN_912; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_946 = 6'h18 == state ? iter_ofm_pre : _GEN_913; // @[control.scala 438:19 194:31]
  wire [31:0] _GEN_947 = 6'h18 == state ? reg_t_4 : _GEN_915; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_948 = 6'h18 == state ? reg_t_5 : _GEN_916; // @[control.scala 438:19 160:37]
  wire  _GEN_949 = 6'h18 == state ? ifm_sel : _GEN_917; // @[control.scala 438:19 379:24]
  wire  _GEN_950 = 6'h18 == state ? resize_load_t : _GEN_918; // @[control.scala 438:19 420:32]
  wire  _GEN_951 = 6'h18 == state ? yolo_finish : _GEN_919; // @[control.scala 438:19 40:28]
  wire  _GEN_952 = 6'h18 == state ? conv_finish : _GEN_920; // @[control.scala 438:19 71:30]
  wire  _GEN_953 = 6'h17 == state ? _T_13 : _GEN_927; // @[control.scala 438:19]
  wire [5:0] _GEN_954 = 6'h17 == state ? {{1'd0}, _GEN_98} : _GEN_926; // @[control.scala 438:19]
  wire [31:0] _GEN_955 = 6'h17 == state ? ifm_addr_fmbase : _GEN_921; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_956 = 6'h17 == state ? ifm_addr_offset : _GEN_922; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_957 = 6'h17 == state ? ifm_send_len : _GEN_923; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_958 = 6'h17 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_924; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_959 = 6'h17 == state ? reg_static : _GEN_925; // @[control.scala 438:19 161:29]
  wire  _GEN_960 = 6'h17 == state ? last_buf_sel : _GEN_928; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_961 = 6'h17 == state ? reg_task : _GEN_929; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_962 = 6'h17 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_930; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_963 = 6'h17 == state ? weight_sel : _GEN_931; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_964 = 6'h17 == state ? wgt_addr_read : _GEN_932; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_965 = 6'h17 == state ? bia_addr_read : _GEN_933; // @[control.scala 438:19 181:32]
  wire  _GEN_966 = 6'h17 == state ? wgt_ddr_read_en : _GEN_934; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_967 = 6'h17 == state ? reg_t_0 : _GEN_935; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_968 = 6'h17 == state ? reg_t_6 : _GEN_936; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_969 = 6'h17 == state ? reg_t_7 : _GEN_937; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_970 = 6'h17 == state ? cnt_t : _GEN_938; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_971 = 6'h17 == state ? pool_cnt : _GEN_939; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_972 = 6'h17 == state ? iter_ifm_post : _GEN_940; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_973 = 6'h17 == state ? iter_div_post : _GEN_941; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_974 = 6'h17 == state ? iter_ofm_post : _GEN_942; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_975 = 6'h17 == state ? iter_ifm_pre : _GEN_943; // @[control.scala 438:19 192:31]
  wire  _GEN_976 = 6'h17 == state ? bottleneck_transfer : _GEN_944; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_977 = 6'h17 == state ? iter_div_pre : _GEN_945; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_978 = 6'h17 == state ? iter_ofm_pre : _GEN_946; // @[control.scala 438:19 194:31]
  wire [31:0] _GEN_979 = 6'h17 == state ? reg_t_4 : _GEN_947; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_980 = 6'h17 == state ? reg_t_5 : _GEN_948; // @[control.scala 438:19 160:37]
  wire  _GEN_981 = 6'h17 == state ? ifm_sel : _GEN_949; // @[control.scala 438:19 379:24]
  wire  _GEN_982 = 6'h17 == state ? resize_load_t : _GEN_950; // @[control.scala 438:19 420:32]
  wire  _GEN_983 = 6'h17 == state ? yolo_finish : _GEN_951; // @[control.scala 438:19 40:28]
  wire  _GEN_984 = 6'h17 == state ? conv_finish : _GEN_952; // @[control.scala 438:19 71:30]
  wire [12:0] _GEN_985 = 6'h16 == state ? _GEN_95 : _GEN_977; // @[control.scala 438:19]
  wire [12:0] _GEN_986 = 6'h16 == state ? _GEN_96 : _GEN_978; // @[control.scala 438:19]
  wire [5:0] _GEN_987 = 6'h16 == state ? 6'h17 : _GEN_954; // @[control.scala 438:19 797:19]
  wire  _GEN_988 = 6'h16 == state ? ifm_send_task_enable : _GEN_953; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_989 = 6'h16 == state ? ifm_addr_fmbase : _GEN_955; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_990 = 6'h16 == state ? ifm_addr_offset : _GEN_956; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_991 = 6'h16 == state ? ifm_send_len : _GEN_957; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_992 = 6'h16 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_958; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_993 = 6'h16 == state ? reg_static : _GEN_959; // @[control.scala 438:19 161:29]
  wire  _GEN_994 = 6'h16 == state ? last_buf_sel : _GEN_960; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_995 = 6'h16 == state ? reg_task : _GEN_961; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_996 = 6'h16 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_962; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_997 = 6'h16 == state ? weight_sel : _GEN_963; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_998 = 6'h16 == state ? wgt_addr_read : _GEN_964; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_999 = 6'h16 == state ? bia_addr_read : _GEN_965; // @[control.scala 438:19 181:32]
  wire  _GEN_1000 = 6'h16 == state ? wgt_ddr_read_en : _GEN_966; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1001 = 6'h16 == state ? reg_t_0 : _GEN_967; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1002 = 6'h16 == state ? reg_t_6 : _GEN_968; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1003 = 6'h16 == state ? reg_t_7 : _GEN_969; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1004 = 6'h16 == state ? cnt_t : _GEN_970; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1005 = 6'h16 == state ? pool_cnt : _GEN_971; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_1006 = 6'h16 == state ? iter_ifm_post : _GEN_972; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1007 = 6'h16 == state ? iter_div_post : _GEN_973; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1008 = 6'h16 == state ? iter_ofm_post : _GEN_974; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1009 = 6'h16 == state ? iter_ifm_pre : _GEN_975; // @[control.scala 438:19 192:31]
  wire  _GEN_1010 = 6'h16 == state ? bottleneck_transfer : _GEN_976; // @[control.scala 438:19 295:38]
  wire [31:0] _GEN_1011 = 6'h16 == state ? reg_t_4 : _GEN_979; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1012 = 6'h16 == state ? reg_t_5 : _GEN_980; // @[control.scala 438:19 160:37]
  wire  _GEN_1013 = 6'h16 == state ? ifm_sel : _GEN_981; // @[control.scala 438:19 379:24]
  wire  _GEN_1014 = 6'h16 == state ? resize_load_t : _GEN_982; // @[control.scala 438:19 420:32]
  wire  _GEN_1015 = 6'h16 == state ? yolo_finish : _GEN_983; // @[control.scala 438:19 40:28]
  wire  _GEN_1016 = 6'h16 == state ? conv_finish : _GEN_984; // @[control.scala 438:19 71:30]
  wire  _GEN_1017 = 6'h15 == state ? bottleneck_en & iter_ifm_pre_t == 13'h1 : _GEN_1010; // @[control.scala 438:19 783:33]
  wire [12:0] _GEN_1018 = 6'h15 == state ? _GEN_92 : _GEN_1009; // @[control.scala 438:19]
  wire [12:0] _GEN_1019 = 6'h15 == state ? _GEN_93 : _GEN_985; // @[control.scala 438:19]
  wire [5:0] _GEN_1020 = 6'h15 == state ? {{1'd0}, _GEN_94} : _GEN_987; // @[control.scala 438:19]
  wire [12:0] _GEN_1021 = 6'h15 == state ? iter_ofm_pre : _GEN_986; // @[control.scala 438:19 194:31]
  wire  _GEN_1022 = 6'h15 == state ? ifm_send_task_enable : _GEN_988; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1023 = 6'h15 == state ? ifm_addr_fmbase : _GEN_989; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1024 = 6'h15 == state ? ifm_addr_offset : _GEN_990; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1025 = 6'h15 == state ? ifm_send_len : _GEN_991; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1026 = 6'h15 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_992; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1027 = 6'h15 == state ? reg_static : _GEN_993; // @[control.scala 438:19 161:29]
  wire  _GEN_1028 = 6'h15 == state ? last_buf_sel : _GEN_994; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1029 = 6'h15 == state ? reg_task : _GEN_995; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1030 = 6'h15 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_996; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1031 = 6'h15 == state ? weight_sel : _GEN_997; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1032 = 6'h15 == state ? wgt_addr_read : _GEN_998; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_1033 = 6'h15 == state ? bia_addr_read : _GEN_999; // @[control.scala 438:19 181:32]
  wire  _GEN_1034 = 6'h15 == state ? wgt_ddr_read_en : _GEN_1000; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1035 = 6'h15 == state ? reg_t_0 : _GEN_1001; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1036 = 6'h15 == state ? reg_t_6 : _GEN_1002; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1037 = 6'h15 == state ? reg_t_7 : _GEN_1003; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1038 = 6'h15 == state ? cnt_t : _GEN_1004; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1039 = 6'h15 == state ? pool_cnt : _GEN_1005; // @[control.scala 438:19 290:27]
  wire [12:0] _GEN_1040 = 6'h15 == state ? iter_ifm_post : _GEN_1006; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1041 = 6'h15 == state ? iter_div_post : _GEN_1007; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1042 = 6'h15 == state ? iter_ofm_post : _GEN_1008; // @[control.scala 438:19 197:32]
  wire [31:0] _GEN_1043 = 6'h15 == state ? reg_t_4 : _GEN_1011; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1044 = 6'h15 == state ? reg_t_5 : _GEN_1012; // @[control.scala 438:19 160:37]
  wire  _GEN_1045 = 6'h15 == state ? ifm_sel : _GEN_1013; // @[control.scala 438:19 379:24]
  wire  _GEN_1046 = 6'h15 == state ? resize_load_t : _GEN_1014; // @[control.scala 438:19 420:32]
  wire  _GEN_1047 = 6'h15 == state ? yolo_finish : _GEN_1015; // @[control.scala 438:19 40:28]
  wire  _GEN_1048 = 6'h15 == state ? conv_finish : _GEN_1016; // @[control.scala 438:19 71:30]
  wire [12:0] _GEN_1049 = 6'h14 == state ? iter_ifm_pre : _GEN_1040; // @[control.scala 438:19 771:27]
  wire [12:0] _GEN_1050 = 6'h14 == state ? iter_div_pre : _GEN_1041; // @[control.scala 438:19 772:27]
  wire [12:0] _GEN_1051 = 6'h14 == state ? iter_ofm_pre : _GEN_1042; // @[control.scala 438:19 773:27]
  wire [5:0] _GEN_1052 = 6'h14 == state ? {{1'd0}, _GEN_90} : _GEN_1020; // @[control.scala 438:19]
  wire [12:0] _GEN_1053 = 6'h14 == state ? _GEN_91 : _GEN_1018; // @[control.scala 438:19]
  wire  _GEN_1054 = 6'h14 == state ? bottleneck_transfer : _GEN_1017; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_1055 = 6'h14 == state ? iter_div_pre : _GEN_1019; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1056 = 6'h14 == state ? iter_ofm_pre : _GEN_1021; // @[control.scala 438:19 194:31]
  wire  _GEN_1057 = 6'h14 == state ? ifm_send_task_enable : _GEN_1022; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1058 = 6'h14 == state ? ifm_addr_fmbase : _GEN_1023; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1059 = 6'h14 == state ? ifm_addr_offset : _GEN_1024; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1060 = 6'h14 == state ? ifm_send_len : _GEN_1025; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1061 = 6'h14 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1026; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1062 = 6'h14 == state ? reg_static : _GEN_1027; // @[control.scala 438:19 161:29]
  wire  _GEN_1063 = 6'h14 == state ? last_buf_sel : _GEN_1028; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1064 = 6'h14 == state ? reg_task : _GEN_1029; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1065 = 6'h14 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1030; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1066 = 6'h14 == state ? weight_sel : _GEN_1031; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1067 = 6'h14 == state ? wgt_addr_read : _GEN_1032; // @[control.scala 438:19 179:32]
  wire [15:0] _GEN_1068 = 6'h14 == state ? bia_addr_read : _GEN_1033; // @[control.scala 438:19 181:32]
  wire  _GEN_1069 = 6'h14 == state ? wgt_ddr_read_en : _GEN_1034; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1070 = 6'h14 == state ? reg_t_0 : _GEN_1035; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1071 = 6'h14 == state ? reg_t_6 : _GEN_1036; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1072 = 6'h14 == state ? reg_t_7 : _GEN_1037; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1073 = 6'h14 == state ? cnt_t : _GEN_1038; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1074 = 6'h14 == state ? pool_cnt : _GEN_1039; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1075 = 6'h14 == state ? reg_t_4 : _GEN_1043; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1076 = 6'h14 == state ? reg_t_5 : _GEN_1044; // @[control.scala 438:19 160:37]
  wire  _GEN_1077 = 6'h14 == state ? ifm_sel : _GEN_1045; // @[control.scala 438:19 379:24]
  wire  _GEN_1078 = 6'h14 == state ? resize_load_t : _GEN_1046; // @[control.scala 438:19 420:32]
  wire  _GEN_1079 = 6'h14 == state ? yolo_finish : _GEN_1047; // @[control.scala 438:19 40:28]
  wire  _GEN_1080 = 6'h14 == state ? conv_finish : _GEN_1048; // @[control.scala 438:19 71:30]
  wire  _GEN_1081 = 6'h13 == state ? _T_67 : wgt_send_task_enable; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1082 = 6'h13 == state ? _GEN_87 : wgt_addr_send; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1083 = 6'h13 == state ? _GEN_88 : _GEN_1067; // @[control.scala 438:19]
  wire [5:0] _GEN_1084 = 6'h13 == state ? _GEN_89 : _GEN_1052; // @[control.scala 438:19]
  wire [12:0] _GEN_1085 = 6'h13 == state ? iter_ifm_post : _GEN_1049; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1086 = 6'h13 == state ? iter_div_post : _GEN_1050; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1087 = 6'h13 == state ? iter_ofm_post : _GEN_1051; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1088 = 6'h13 == state ? iter_ifm_pre : _GEN_1053; // @[control.scala 438:19 192:31]
  wire  _GEN_1089 = 6'h13 == state ? bottleneck_transfer : _GEN_1054; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_1090 = 6'h13 == state ? iter_div_pre : _GEN_1055; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1091 = 6'h13 == state ? iter_ofm_pre : _GEN_1056; // @[control.scala 438:19 194:31]
  wire  _GEN_1092 = 6'h13 == state ? ifm_send_task_enable : _GEN_1057; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1093 = 6'h13 == state ? ifm_addr_fmbase : _GEN_1058; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1094 = 6'h13 == state ? ifm_addr_offset : _GEN_1059; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1095 = 6'h13 == state ? ifm_send_len : _GEN_1060; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1096 = 6'h13 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1061; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1097 = 6'h13 == state ? reg_static : _GEN_1062; // @[control.scala 438:19 161:29]
  wire  _GEN_1098 = 6'h13 == state ? last_buf_sel : _GEN_1063; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1099 = 6'h13 == state ? reg_task : _GEN_1064; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1100 = 6'h13 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1065; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1101 = 6'h13 == state ? weight_sel : _GEN_1066; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1102 = 6'h13 == state ? bia_addr_read : _GEN_1068; // @[control.scala 438:19 181:32]
  wire  _GEN_1103 = 6'h13 == state ? wgt_ddr_read_en : _GEN_1069; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1104 = 6'h13 == state ? reg_t_0 : _GEN_1070; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1105 = 6'h13 == state ? reg_t_6 : _GEN_1071; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1106 = 6'h13 == state ? reg_t_7 : _GEN_1072; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1107 = 6'h13 == state ? cnt_t : _GEN_1073; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1108 = 6'h13 == state ? pool_cnt : _GEN_1074; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1109 = 6'h13 == state ? reg_t_4 : _GEN_1075; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1110 = 6'h13 == state ? reg_t_5 : _GEN_1076; // @[control.scala 438:19 160:37]
  wire  _GEN_1111 = 6'h13 == state ? ifm_sel : _GEN_1077; // @[control.scala 438:19 379:24]
  wire  _GEN_1112 = 6'h13 == state ? resize_load_t : _GEN_1078; // @[control.scala 438:19 420:32]
  wire  _GEN_1113 = 6'h13 == state ? yolo_finish : _GEN_1079; // @[control.scala 438:19 40:28]
  wire  _GEN_1114 = 6'h13 == state ? conv_finish : _GEN_1080; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_1115 = 6'h12 == state ? 6'h13 : _GEN_1084; // @[control.scala 438:19 744:19]
  wire [31:0] _GEN_1116 = 6'h12 == state ? _GEN_84 : ofm_addr_offset; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1117 = 6'h12 == state ? {{13'd0}, _GEN_85} : ofm_recv_len; // @[control.scala 438:19 367:31]
  wire  _GEN_1118 = 6'h12 == state ? wgt_send_task_enable : _GEN_1081; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1119 = 6'h12 == state ? wgt_addr_send : _GEN_1082; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1120 = 6'h12 == state ? wgt_addr_read : _GEN_1083; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1121 = 6'h12 == state ? iter_ifm_post : _GEN_1085; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1122 = 6'h12 == state ? iter_div_post : _GEN_1086; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1123 = 6'h12 == state ? iter_ofm_post : _GEN_1087; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1124 = 6'h12 == state ? iter_ifm_pre : _GEN_1088; // @[control.scala 438:19 192:31]
  wire  _GEN_1125 = 6'h12 == state ? bottleneck_transfer : _GEN_1089; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_1126 = 6'h12 == state ? iter_div_pre : _GEN_1090; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1127 = 6'h12 == state ? iter_ofm_pre : _GEN_1091; // @[control.scala 438:19 194:31]
  wire  _GEN_1128 = 6'h12 == state ? ifm_send_task_enable : _GEN_1092; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1129 = 6'h12 == state ? ifm_addr_fmbase : _GEN_1093; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1130 = 6'h12 == state ? ifm_addr_offset : _GEN_1094; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1131 = 6'h12 == state ? ifm_send_len : _GEN_1095; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1132 = 6'h12 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1096; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1133 = 6'h12 == state ? reg_static : _GEN_1097; // @[control.scala 438:19 161:29]
  wire  _GEN_1134 = 6'h12 == state ? last_buf_sel : _GEN_1098; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1135 = 6'h12 == state ? reg_task : _GEN_1099; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1136 = 6'h12 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1100; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1137 = 6'h12 == state ? weight_sel : _GEN_1101; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1138 = 6'h12 == state ? bia_addr_read : _GEN_1102; // @[control.scala 438:19 181:32]
  wire  _GEN_1139 = 6'h12 == state ? wgt_ddr_read_en : _GEN_1103; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1140 = 6'h12 == state ? reg_t_0 : _GEN_1104; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1141 = 6'h12 == state ? reg_t_6 : _GEN_1105; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1142 = 6'h12 == state ? reg_t_7 : _GEN_1106; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1143 = 6'h12 == state ? cnt_t : _GEN_1107; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1144 = 6'h12 == state ? pool_cnt : _GEN_1108; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1145 = 6'h12 == state ? reg_t_4 : _GEN_1109; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1146 = 6'h12 == state ? reg_t_5 : _GEN_1110; // @[control.scala 438:19 160:37]
  wire  _GEN_1147 = 6'h12 == state ? ifm_sel : _GEN_1111; // @[control.scala 438:19 379:24]
  wire  _GEN_1148 = 6'h12 == state ? resize_load_t : _GEN_1112; // @[control.scala 438:19 420:32]
  wire  _GEN_1149 = 6'h12 == state ? yolo_finish : _GEN_1113; // @[control.scala 438:19 40:28]
  wire  _GEN_1150 = 6'h12 == state ? conv_finish : _GEN_1114; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1151 = 6'h11 == state ? _ofm_addr_fmbase_T : ofm_addr_fmbase; // @[control.scala 438:19 733:29 365:34]
  wire [31:0] _GEN_1152 = 6'h11 == state ? _GEN_81 : _GEN_1116; // @[control.scala 438:19]
  wire [31:0] _GEN_1153 = 6'h11 == state ? _GEN_82 : _GEN_1117; // @[control.scala 438:19]
  wire [5:0] _GEN_1154 = 6'h11 == state ? {{1'd0}, _GEN_83} : _GEN_1115; // @[control.scala 438:19]
  wire  _GEN_1155 = 6'h11 == state ? wgt_send_task_enable : _GEN_1118; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1156 = 6'h11 == state ? wgt_addr_send : _GEN_1119; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1157 = 6'h11 == state ? wgt_addr_read : _GEN_1120; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1158 = 6'h11 == state ? iter_ifm_post : _GEN_1121; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1159 = 6'h11 == state ? iter_div_post : _GEN_1122; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1160 = 6'h11 == state ? iter_ofm_post : _GEN_1123; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1161 = 6'h11 == state ? iter_ifm_pre : _GEN_1124; // @[control.scala 438:19 192:31]
  wire  _GEN_1162 = 6'h11 == state ? bottleneck_transfer : _GEN_1125; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_1163 = 6'h11 == state ? iter_div_pre : _GEN_1126; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1164 = 6'h11 == state ? iter_ofm_pre : _GEN_1127; // @[control.scala 438:19 194:31]
  wire  _GEN_1165 = 6'h11 == state ? ifm_send_task_enable : _GEN_1128; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1166 = 6'h11 == state ? ifm_addr_fmbase : _GEN_1129; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1167 = 6'h11 == state ? ifm_addr_offset : _GEN_1130; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1168 = 6'h11 == state ? ifm_send_len : _GEN_1131; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1169 = 6'h11 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1132; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1170 = 6'h11 == state ? reg_static : _GEN_1133; // @[control.scala 438:19 161:29]
  wire  _GEN_1171 = 6'h11 == state ? last_buf_sel : _GEN_1134; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1172 = 6'h11 == state ? reg_task : _GEN_1135; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1173 = 6'h11 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1136; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1174 = 6'h11 == state ? weight_sel : _GEN_1137; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1175 = 6'h11 == state ? bia_addr_read : _GEN_1138; // @[control.scala 438:19 181:32]
  wire  _GEN_1176 = 6'h11 == state ? wgt_ddr_read_en : _GEN_1139; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1177 = 6'h11 == state ? reg_t_0 : _GEN_1140; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1178 = 6'h11 == state ? reg_t_6 : _GEN_1141; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1179 = 6'h11 == state ? reg_t_7 : _GEN_1142; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1180 = 6'h11 == state ? cnt_t : _GEN_1143; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1181 = 6'h11 == state ? pool_cnt : _GEN_1144; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1182 = 6'h11 == state ? reg_t_4 : _GEN_1145; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1183 = 6'h11 == state ? reg_t_5 : _GEN_1146; // @[control.scala 438:19 160:37]
  wire  _GEN_1184 = 6'h11 == state ? ifm_sel : _GEN_1147; // @[control.scala 438:19 379:24]
  wire  _GEN_1185 = 6'h11 == state ? resize_load_t : _GEN_1148; // @[control.scala 438:19 420:32]
  wire  _GEN_1186 = 6'h11 == state ? yolo_finish : _GEN_1149; // @[control.scala 438:19 40:28]
  wire  _GEN_1187 = 6'h11 == state ? conv_finish : _GEN_1150; // @[control.scala 438:19 71:30]
  wire  _GEN_1188 = 6'h10 == state ? _T_58 : ofm_recv_task_enable; // @[control.scala 438:19 358:39]
  wire [5:0] _GEN_1189 = 6'h10 == state ? {{1'd0}, _GEN_79} : _GEN_1154; // @[control.scala 438:19]
  wire  _GEN_1190 = 6'h10 == state ? _GEN_80 : first_ofm_recv_stop; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1191 = 6'h10 == state ? ofm_addr_fmbase : _GEN_1151; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1192 = 6'h10 == state ? ofm_addr_offset : _GEN_1152; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1193 = 6'h10 == state ? ofm_recv_len : _GEN_1153; // @[control.scala 438:19 367:31]
  wire  _GEN_1194 = 6'h10 == state ? wgt_send_task_enable : _GEN_1155; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1195 = 6'h10 == state ? wgt_addr_send : _GEN_1156; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1196 = 6'h10 == state ? wgt_addr_read : _GEN_1157; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1197 = 6'h10 == state ? iter_ifm_post : _GEN_1158; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1198 = 6'h10 == state ? iter_div_post : _GEN_1159; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1199 = 6'h10 == state ? iter_ofm_post : _GEN_1160; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1200 = 6'h10 == state ? iter_ifm_pre : _GEN_1161; // @[control.scala 438:19 192:31]
  wire  _GEN_1201 = 6'h10 == state ? bottleneck_transfer : _GEN_1162; // @[control.scala 438:19 295:38]
  wire [12:0] _GEN_1202 = 6'h10 == state ? iter_div_pre : _GEN_1163; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1203 = 6'h10 == state ? iter_ofm_pre : _GEN_1164; // @[control.scala 438:19 194:31]
  wire  _GEN_1204 = 6'h10 == state ? ifm_send_task_enable : _GEN_1165; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1205 = 6'h10 == state ? ifm_addr_fmbase : _GEN_1166; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1206 = 6'h10 == state ? ifm_addr_offset : _GEN_1167; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1207 = 6'h10 == state ? ifm_send_len : _GEN_1168; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1208 = 6'h10 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1169; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1209 = 6'h10 == state ? reg_static : _GEN_1170; // @[control.scala 438:19 161:29]
  wire  _GEN_1210 = 6'h10 == state ? last_buf_sel : _GEN_1171; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1211 = 6'h10 == state ? reg_task : _GEN_1172; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1212 = 6'h10 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1173; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1213 = 6'h10 == state ? weight_sel : _GEN_1174; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1214 = 6'h10 == state ? bia_addr_read : _GEN_1175; // @[control.scala 438:19 181:32]
  wire  _GEN_1215 = 6'h10 == state ? wgt_ddr_read_en : _GEN_1176; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1216 = 6'h10 == state ? reg_t_0 : _GEN_1177; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1217 = 6'h10 == state ? reg_t_6 : _GEN_1178; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1218 = 6'h10 == state ? reg_t_7 : _GEN_1179; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1219 = 6'h10 == state ? cnt_t : _GEN_1180; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1220 = 6'h10 == state ? pool_cnt : _GEN_1181; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1221 = 6'h10 == state ? reg_t_4 : _GEN_1182; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1222 = 6'h10 == state ? reg_t_5 : _GEN_1183; // @[control.scala 438:19 160:37]
  wire  _GEN_1223 = 6'h10 == state ? ifm_sel : _GEN_1184; // @[control.scala 438:19 379:24]
  wire  _GEN_1224 = 6'h10 == state ? resize_load_t : _GEN_1185; // @[control.scala 438:19 420:32]
  wire  _GEN_1225 = 6'h10 == state ? yolo_finish : _GEN_1186; // @[control.scala 438:19 40:28]
  wire  _GEN_1226 = 6'h10 == state ? conv_finish : _GEN_1187; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_1227 = 6'hf == state ? {{1'd0}, _GEN_75} : _GEN_1189; // @[control.scala 438:19]
  wire  _GEN_1228 = 6'hf == state ? _GEN_76 : _GEN_1201; // @[control.scala 438:19]
  wire  _GEN_1229 = 6'hf == state ? _GEN_77 : bottleneck_ready; // @[control.scala 438:19 296:35]
  wire  _GEN_1230 = 6'hf == state ? ofm_recv_task_enable : _GEN_1188; // @[control.scala 438:19 358:39]
  wire  _GEN_1231 = 6'hf == state ? first_ofm_recv_stop : _GEN_1190; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1232 = 6'hf == state ? ofm_addr_fmbase : _GEN_1191; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1233 = 6'hf == state ? ofm_addr_offset : _GEN_1192; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1234 = 6'hf == state ? ofm_recv_len : _GEN_1193; // @[control.scala 438:19 367:31]
  wire  _GEN_1235 = 6'hf == state ? wgt_send_task_enable : _GEN_1194; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1236 = 6'hf == state ? wgt_addr_send : _GEN_1195; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1237 = 6'hf == state ? wgt_addr_read : _GEN_1196; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1238 = 6'hf == state ? iter_ifm_post : _GEN_1197; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1239 = 6'hf == state ? iter_div_post : _GEN_1198; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1240 = 6'hf == state ? iter_ofm_post : _GEN_1199; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1241 = 6'hf == state ? iter_ifm_pre : _GEN_1200; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1242 = 6'hf == state ? iter_div_pre : _GEN_1202; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1243 = 6'hf == state ? iter_ofm_pre : _GEN_1203; // @[control.scala 438:19 194:31]
  wire  _GEN_1244 = 6'hf == state ? ifm_send_task_enable : _GEN_1204; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1245 = 6'hf == state ? ifm_addr_fmbase : _GEN_1205; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1246 = 6'hf == state ? ifm_addr_offset : _GEN_1206; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1247 = 6'hf == state ? ifm_send_len : _GEN_1207; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1248 = 6'hf == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1208; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1249 = 6'hf == state ? reg_static : _GEN_1209; // @[control.scala 438:19 161:29]
  wire  _GEN_1250 = 6'hf == state ? last_buf_sel : _GEN_1210; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1251 = 6'hf == state ? reg_task : _GEN_1211; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1252 = 6'hf == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1212; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1253 = 6'hf == state ? weight_sel : _GEN_1213; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1254 = 6'hf == state ? bia_addr_read : _GEN_1214; // @[control.scala 438:19 181:32]
  wire  _GEN_1255 = 6'hf == state ? wgt_ddr_read_en : _GEN_1215; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1256 = 6'hf == state ? reg_t_0 : _GEN_1216; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1257 = 6'hf == state ? reg_t_6 : _GEN_1217; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1258 = 6'hf == state ? reg_t_7 : _GEN_1218; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1259 = 6'hf == state ? cnt_t : _GEN_1219; // @[control.scala 438:19 163:24]
  wire [1:0] _GEN_1260 = 6'hf == state ? pool_cnt : _GEN_1220; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1261 = 6'hf == state ? reg_t_4 : _GEN_1221; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1262 = 6'hf == state ? reg_t_5 : _GEN_1222; // @[control.scala 438:19 160:37]
  wire  _GEN_1263 = 6'hf == state ? ifm_sel : _GEN_1223; // @[control.scala 438:19 379:24]
  wire  _GEN_1264 = 6'hf == state ? resize_load_t : _GEN_1224; // @[control.scala 438:19 420:32]
  wire  _GEN_1265 = 6'hf == state ? yolo_finish : _GEN_1225; // @[control.scala 438:19 40:28]
  wire  _GEN_1266 = 6'hf == state ? conv_finish : _GEN_1226; // @[control.scala 438:19 71:30]
  wire [4:0] _GEN_1267 = 6'he == state ? _GEN_2 : _GEN_1259; // @[control.scala 438:19]
  wire [5:0] _GEN_1268 = 6'he == state ? _GEN_70 : _GEN_1227; // @[control.scala 438:19]
  wire [31:0] _GEN_1269 = 6'he == state ? _GEN_71 : _GEN_1256; // @[control.scala 438:19]
  wire  _GEN_1270 = 6'he == state ? bottleneck_transfer : _GEN_1228; // @[control.scala 438:19 295:38]
  wire  _GEN_1271 = 6'he == state ? bottleneck_ready : _GEN_1229; // @[control.scala 438:19 296:35]
  wire  _GEN_1272 = 6'he == state ? ofm_recv_task_enable : _GEN_1230; // @[control.scala 438:19 358:39]
  wire  _GEN_1273 = 6'he == state ? first_ofm_recv_stop : _GEN_1231; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1274 = 6'he == state ? ofm_addr_fmbase : _GEN_1232; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1275 = 6'he == state ? ofm_addr_offset : _GEN_1233; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1276 = 6'he == state ? ofm_recv_len : _GEN_1234; // @[control.scala 438:19 367:31]
  wire  _GEN_1277 = 6'he == state ? wgt_send_task_enable : _GEN_1235; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1278 = 6'he == state ? wgt_addr_send : _GEN_1236; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1279 = 6'he == state ? wgt_addr_read : _GEN_1237; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1280 = 6'he == state ? iter_ifm_post : _GEN_1238; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1281 = 6'he == state ? iter_div_post : _GEN_1239; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1282 = 6'he == state ? iter_ofm_post : _GEN_1240; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1283 = 6'he == state ? iter_ifm_pre : _GEN_1241; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1284 = 6'he == state ? iter_div_pre : _GEN_1242; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1285 = 6'he == state ? iter_ofm_pre : _GEN_1243; // @[control.scala 438:19 194:31]
  wire  _GEN_1286 = 6'he == state ? ifm_send_task_enable : _GEN_1244; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1287 = 6'he == state ? ifm_addr_fmbase : _GEN_1245; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1288 = 6'he == state ? ifm_addr_offset : _GEN_1246; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1289 = 6'he == state ? ifm_send_len : _GEN_1247; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1290 = 6'he == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1248; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1291 = 6'he == state ? reg_static : _GEN_1249; // @[control.scala 438:19 161:29]
  wire  _GEN_1292 = 6'he == state ? last_buf_sel : _GEN_1250; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1293 = 6'he == state ? reg_task : _GEN_1251; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1294 = 6'he == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1252; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1295 = 6'he == state ? weight_sel : _GEN_1253; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1296 = 6'he == state ? bia_addr_read : _GEN_1254; // @[control.scala 438:19 181:32]
  wire  _GEN_1297 = 6'he == state ? wgt_ddr_read_en : _GEN_1255; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1298 = 6'he == state ? reg_t_6 : _GEN_1257; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1299 = 6'he == state ? reg_t_7 : _GEN_1258; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1300 = 6'he == state ? pool_cnt : _GEN_1260; // @[control.scala 438:19 290:27]
  wire [31:0] _GEN_1301 = 6'he == state ? reg_t_4 : _GEN_1261; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1302 = 6'he == state ? reg_t_5 : _GEN_1262; // @[control.scala 438:19 160:37]
  wire  _GEN_1303 = 6'he == state ? ifm_sel : _GEN_1263; // @[control.scala 438:19 379:24]
  wire  _GEN_1304 = 6'he == state ? resize_load_t : _GEN_1264; // @[control.scala 438:19 420:32]
  wire  _GEN_1305 = 6'he == state ? yolo_finish : _GEN_1265; // @[control.scala 438:19 40:28]
  wire  _GEN_1306 = 6'he == state ? conv_finish : _GEN_1266; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1307 = 6'hd == state ? _GEN_67 : _GEN_1301; // @[control.scala 438:19]
  wire [31:0] _GEN_1308 = 6'hd == state ? _GEN_68 : _GEN_1302; // @[control.scala 438:19]
  wire [31:0] _GEN_1309 = 6'hd == state ? _reg_t_3_T_2 : reg_t_3; // @[control.scala 438:19 689:22 160:37]
  wire [31:0] _GEN_1310 = 6'hd == state ? _reg_t_0_T_4 : _GEN_1269; // @[control.scala 438:19 690:22]
  wire [4:0] _GEN_1311 = 6'hd == state ? 5'h0 : _GEN_1267; // @[control.scala 438:19 691:19]
  wire [5:0] _GEN_1312 = 6'hd == state ? 6'he : _GEN_1268; // @[control.scala 438:19 692:19]
  wire  _GEN_1313 = 6'hd == state ? bottleneck_transfer : _GEN_1270; // @[control.scala 438:19 295:38]
  wire  _GEN_1314 = 6'hd == state ? bottleneck_ready : _GEN_1271; // @[control.scala 438:19 296:35]
  wire  _GEN_1315 = 6'hd == state ? ofm_recv_task_enable : _GEN_1272; // @[control.scala 438:19 358:39]
  wire  _GEN_1316 = 6'hd == state ? first_ofm_recv_stop : _GEN_1273; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1317 = 6'hd == state ? ofm_addr_fmbase : _GEN_1274; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1318 = 6'hd == state ? ofm_addr_offset : _GEN_1275; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1319 = 6'hd == state ? ofm_recv_len : _GEN_1276; // @[control.scala 438:19 367:31]
  wire  _GEN_1320 = 6'hd == state ? wgt_send_task_enable : _GEN_1277; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1321 = 6'hd == state ? wgt_addr_send : _GEN_1278; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1322 = 6'hd == state ? wgt_addr_read : _GEN_1279; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1323 = 6'hd == state ? iter_ifm_post : _GEN_1280; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1324 = 6'hd == state ? iter_div_post : _GEN_1281; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1325 = 6'hd == state ? iter_ofm_post : _GEN_1282; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1326 = 6'hd == state ? iter_ifm_pre : _GEN_1283; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1327 = 6'hd == state ? iter_div_pre : _GEN_1284; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1328 = 6'hd == state ? iter_ofm_pre : _GEN_1285; // @[control.scala 438:19 194:31]
  wire  _GEN_1329 = 6'hd == state ? ifm_send_task_enable : _GEN_1286; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1330 = 6'hd == state ? ifm_addr_fmbase : _GEN_1287; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1331 = 6'hd == state ? ifm_addr_offset : _GEN_1288; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1332 = 6'hd == state ? ifm_send_len : _GEN_1289; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1333 = 6'hd == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1290; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1334 = 6'hd == state ? reg_static : _GEN_1291; // @[control.scala 438:19 161:29]
  wire  _GEN_1335 = 6'hd == state ? last_buf_sel : _GEN_1292; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1336 = 6'hd == state ? reg_task : _GEN_1293; // @[control.scala 438:19 162:27]
  wire [25:0] _GEN_1337 = 6'hd == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1294; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1338 = 6'hd == state ? weight_sel : _GEN_1295; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1339 = 6'hd == state ? bia_addr_read : _GEN_1296; // @[control.scala 438:19 181:32]
  wire  _GEN_1340 = 6'hd == state ? wgt_ddr_read_en : _GEN_1297; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1341 = 6'hd == state ? reg_t_6 : _GEN_1298; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1342 = 6'hd == state ? reg_t_7 : _GEN_1299; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1343 = 6'hd == state ? pool_cnt : _GEN_1300; // @[control.scala 438:19 290:27]
  wire  _GEN_1344 = 6'hd == state ? ifm_sel : _GEN_1303; // @[control.scala 438:19 379:24]
  wire  _GEN_1345 = 6'hd == state ? resize_load_t : _GEN_1304; // @[control.scala 438:19 420:32]
  wire  _GEN_1346 = 6'hd == state ? yolo_finish : _GEN_1305; // @[control.scala 438:19 40:28]
  wire  _GEN_1347 = 6'hd == state ? conv_finish : _GEN_1306; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1348 = 6'hc == state ? _GEN_62 : _GEN_1334; // @[control.scala 438:19]
  wire [31:0] _GEN_1349 = 6'hc == state ? {{12'd0}, _GEN_66} : _GEN_1336; // @[control.scala 438:19]
  wire [5:0] _GEN_1350 = 6'hc == state ? 6'hd : _GEN_1312; // @[control.scala 438:19 677:19]
  wire [31:0] _GEN_1351 = 6'hc == state ? reg_t_4 : _GEN_1307; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1352 = 6'hc == state ? reg_t_5 : _GEN_1308; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1353 = 6'hc == state ? reg_t_3 : _GEN_1309; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1354 = 6'hc == state ? reg_t_0 : _GEN_1310; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1355 = 6'hc == state ? cnt_t : _GEN_1311; // @[control.scala 438:19 163:24]
  wire  _GEN_1356 = 6'hc == state ? bottleneck_transfer : _GEN_1313; // @[control.scala 438:19 295:38]
  wire  _GEN_1357 = 6'hc == state ? bottleneck_ready : _GEN_1314; // @[control.scala 438:19 296:35]
  wire  _GEN_1358 = 6'hc == state ? ofm_recv_task_enable : _GEN_1315; // @[control.scala 438:19 358:39]
  wire  _GEN_1359 = 6'hc == state ? first_ofm_recv_stop : _GEN_1316; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1360 = 6'hc == state ? ofm_addr_fmbase : _GEN_1317; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1361 = 6'hc == state ? ofm_addr_offset : _GEN_1318; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1362 = 6'hc == state ? ofm_recv_len : _GEN_1319; // @[control.scala 438:19 367:31]
  wire  _GEN_1363 = 6'hc == state ? wgt_send_task_enable : _GEN_1320; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1364 = 6'hc == state ? wgt_addr_send : _GEN_1321; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1365 = 6'hc == state ? wgt_addr_read : _GEN_1322; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1366 = 6'hc == state ? iter_ifm_post : _GEN_1323; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1367 = 6'hc == state ? iter_div_post : _GEN_1324; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1368 = 6'hc == state ? iter_ofm_post : _GEN_1325; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1369 = 6'hc == state ? iter_ifm_pre : _GEN_1326; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1370 = 6'hc == state ? iter_div_pre : _GEN_1327; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1371 = 6'hc == state ? iter_ofm_pre : _GEN_1328; // @[control.scala 438:19 194:31]
  wire  _GEN_1372 = 6'hc == state ? ifm_send_task_enable : _GEN_1329; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1373 = 6'hc == state ? ifm_addr_fmbase : _GEN_1330; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1374 = 6'hc == state ? ifm_addr_offset : _GEN_1331; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1375 = 6'hc == state ? ifm_send_len : _GEN_1332; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1376 = 6'hc == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1333; // @[control.scala 438:19 425:46]
  wire  _GEN_1377 = 6'hc == state ? last_buf_sel : _GEN_1335; // @[control.scala 438:19 182:31]
  wire [25:0] _GEN_1378 = 6'hc == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1337; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1379 = 6'hc == state ? weight_sel : _GEN_1338; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1380 = 6'hc == state ? bia_addr_read : _GEN_1339; // @[control.scala 438:19 181:32]
  wire  _GEN_1381 = 6'hc == state ? wgt_ddr_read_en : _GEN_1340; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1382 = 6'hc == state ? reg_t_6 : _GEN_1341; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1383 = 6'hc == state ? reg_t_7 : _GEN_1342; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1384 = 6'hc == state ? pool_cnt : _GEN_1343; // @[control.scala 438:19 290:27]
  wire  _GEN_1385 = 6'hc == state ? ifm_sel : _GEN_1344; // @[control.scala 438:19 379:24]
  wire  _GEN_1386 = 6'hc == state ? resize_load_t : _GEN_1345; // @[control.scala 438:19 420:32]
  wire  _GEN_1387 = 6'hc == state ? yolo_finish : _GEN_1346; // @[control.scala 438:19 40:28]
  wire  _GEN_1388 = 6'hc == state ? conv_finish : _GEN_1347; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1389 = 6'hb == state ? _GEN_55 : _GEN_1348; // @[control.scala 438:19]
  wire [5:0] _GEN_1390 = 6'hb == state ? 6'hc : _GEN_1350; // @[control.scala 438:19 630:18]
  wire [31:0] _GEN_1391 = 6'hb == state ? reg_task : _GEN_1349; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1392 = 6'hb == state ? reg_t_4 : _GEN_1351; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1393 = 6'hb == state ? reg_t_5 : _GEN_1352; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1394 = 6'hb == state ? reg_t_3 : _GEN_1353; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1395 = 6'hb == state ? reg_t_0 : _GEN_1354; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1396 = 6'hb == state ? cnt_t : _GEN_1355; // @[control.scala 438:19 163:24]
  wire  _GEN_1397 = 6'hb == state ? bottleneck_transfer : _GEN_1356; // @[control.scala 438:19 295:38]
  wire  _GEN_1398 = 6'hb == state ? bottleneck_ready : _GEN_1357; // @[control.scala 438:19 296:35]
  wire  _GEN_1399 = 6'hb == state ? ofm_recv_task_enable : _GEN_1358; // @[control.scala 438:19 358:39]
  wire  _GEN_1400 = 6'hb == state ? first_ofm_recv_stop : _GEN_1359; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1401 = 6'hb == state ? ofm_addr_fmbase : _GEN_1360; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1402 = 6'hb == state ? ofm_addr_offset : _GEN_1361; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1403 = 6'hb == state ? ofm_recv_len : _GEN_1362; // @[control.scala 438:19 367:31]
  wire  _GEN_1404 = 6'hb == state ? wgt_send_task_enable : _GEN_1363; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1405 = 6'hb == state ? wgt_addr_send : _GEN_1364; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1406 = 6'hb == state ? wgt_addr_read : _GEN_1365; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1407 = 6'hb == state ? iter_ifm_post : _GEN_1366; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1408 = 6'hb == state ? iter_div_post : _GEN_1367; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1409 = 6'hb == state ? iter_ofm_post : _GEN_1368; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1410 = 6'hb == state ? iter_ifm_pre : _GEN_1369; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1411 = 6'hb == state ? iter_div_pre : _GEN_1370; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1412 = 6'hb == state ? iter_ofm_pre : _GEN_1371; // @[control.scala 438:19 194:31]
  wire  _GEN_1413 = 6'hb == state ? ifm_send_task_enable : _GEN_1372; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1414 = 6'hb == state ? ifm_addr_fmbase : _GEN_1373; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1415 = 6'hb == state ? ifm_addr_offset : _GEN_1374; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1416 = 6'hb == state ? ifm_send_len : _GEN_1375; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1417 = 6'hb == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1376; // @[control.scala 438:19 425:46]
  wire  _GEN_1418 = 6'hb == state ? last_buf_sel : _GEN_1377; // @[control.scala 438:19 182:31]
  wire [25:0] _GEN_1419 = 6'hb == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1378; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1420 = 6'hb == state ? weight_sel : _GEN_1379; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1421 = 6'hb == state ? bia_addr_read : _GEN_1380; // @[control.scala 438:19 181:32]
  wire  _GEN_1422 = 6'hb == state ? wgt_ddr_read_en : _GEN_1381; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1423 = 6'hb == state ? reg_t_6 : _GEN_1382; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1424 = 6'hb == state ? reg_t_7 : _GEN_1383; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1425 = 6'hb == state ? pool_cnt : _GEN_1384; // @[control.scala 438:19 290:27]
  wire  _GEN_1426 = 6'hb == state ? ifm_sel : _GEN_1385; // @[control.scala 438:19 379:24]
  wire  _GEN_1427 = 6'hb == state ? resize_load_t : _GEN_1386; // @[control.scala 438:19 420:32]
  wire  _GEN_1428 = 6'hb == state ? yolo_finish : _GEN_1387; // @[control.scala 438:19 40:28]
  wire  _GEN_1429 = 6'hb == state ? conv_finish : _GEN_1388; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1430 = 6'ha == state ? _GEN_52 : _GEN_1389; // @[control.scala 438:19]
  wire  _GEN_1431 = 6'ha == state ? _T_28 : _GEN_1418; // @[control.scala 438:19 619:26]
  wire [5:0] _GEN_1432 = 6'ha == state ? 6'hb : _GEN_1390; // @[control.scala 438:19 620:19]
  wire [31:0] _GEN_1433 = 6'ha == state ? reg_task : _GEN_1391; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1434 = 6'ha == state ? reg_t_4 : _GEN_1392; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1435 = 6'ha == state ? reg_t_5 : _GEN_1393; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1436 = 6'ha == state ? reg_t_3 : _GEN_1394; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1437 = 6'ha == state ? reg_t_0 : _GEN_1395; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1438 = 6'ha == state ? cnt_t : _GEN_1396; // @[control.scala 438:19 163:24]
  wire  _GEN_1439 = 6'ha == state ? bottleneck_transfer : _GEN_1397; // @[control.scala 438:19 295:38]
  wire  _GEN_1440 = 6'ha == state ? bottleneck_ready : _GEN_1398; // @[control.scala 438:19 296:35]
  wire  _GEN_1441 = 6'ha == state ? ofm_recv_task_enable : _GEN_1399; // @[control.scala 438:19 358:39]
  wire  _GEN_1442 = 6'ha == state ? first_ofm_recv_stop : _GEN_1400; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1443 = 6'ha == state ? ofm_addr_fmbase : _GEN_1401; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1444 = 6'ha == state ? ofm_addr_offset : _GEN_1402; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1445 = 6'ha == state ? ofm_recv_len : _GEN_1403; // @[control.scala 438:19 367:31]
  wire  _GEN_1446 = 6'ha == state ? wgt_send_task_enable : _GEN_1404; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1447 = 6'ha == state ? wgt_addr_send : _GEN_1405; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1448 = 6'ha == state ? wgt_addr_read : _GEN_1406; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1449 = 6'ha == state ? iter_ifm_post : _GEN_1407; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1450 = 6'ha == state ? iter_div_post : _GEN_1408; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1451 = 6'ha == state ? iter_ofm_post : _GEN_1409; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1452 = 6'ha == state ? iter_ifm_pre : _GEN_1410; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1453 = 6'ha == state ? iter_div_pre : _GEN_1411; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1454 = 6'ha == state ? iter_ofm_pre : _GEN_1412; // @[control.scala 438:19 194:31]
  wire  _GEN_1455 = 6'ha == state ? ifm_send_task_enable : _GEN_1413; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1456 = 6'ha == state ? ifm_addr_fmbase : _GEN_1414; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1457 = 6'ha == state ? ifm_addr_offset : _GEN_1415; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1458 = 6'ha == state ? ifm_send_len : _GEN_1416; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1459 = 6'ha == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1417; // @[control.scala 438:19 425:46]
  wire [25:0] _GEN_1460 = 6'ha == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1419; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1461 = 6'ha == state ? weight_sel : _GEN_1420; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1462 = 6'ha == state ? bia_addr_read : _GEN_1421; // @[control.scala 438:19 181:32]
  wire  _GEN_1463 = 6'ha == state ? wgt_ddr_read_en : _GEN_1422; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1464 = 6'ha == state ? reg_t_6 : _GEN_1423; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1465 = 6'ha == state ? reg_t_7 : _GEN_1424; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1466 = 6'ha == state ? pool_cnt : _GEN_1425; // @[control.scala 438:19 290:27]
  wire  _GEN_1467 = 6'ha == state ? ifm_sel : _GEN_1426; // @[control.scala 438:19 379:24]
  wire  _GEN_1468 = 6'ha == state ? resize_load_t : _GEN_1427; // @[control.scala 438:19 420:32]
  wire  _GEN_1469 = 6'ha == state ? yolo_finish : _GEN_1428; // @[control.scala 438:19 40:28]
  wire  _GEN_1470 = 6'ha == state ? conv_finish : _GEN_1429; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1471 = 6'h9 == state ? _GEN_51 : _GEN_1430; // @[control.scala 438:19]
  wire [5:0] _GEN_1472 = 6'h9 == state ? 6'ha : _GEN_1432; // @[control.scala 438:19 613:19]
  wire  _GEN_1473 = 6'h9 == state ? last_buf_sel : _GEN_1431; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1474 = 6'h9 == state ? reg_task : _GEN_1433; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1475 = 6'h9 == state ? reg_t_4 : _GEN_1434; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1476 = 6'h9 == state ? reg_t_5 : _GEN_1435; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1477 = 6'h9 == state ? reg_t_3 : _GEN_1436; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1478 = 6'h9 == state ? reg_t_0 : _GEN_1437; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1479 = 6'h9 == state ? cnt_t : _GEN_1438; // @[control.scala 438:19 163:24]
  wire  _GEN_1480 = 6'h9 == state ? bottleneck_transfer : _GEN_1439; // @[control.scala 438:19 295:38]
  wire  _GEN_1481 = 6'h9 == state ? bottleneck_ready : _GEN_1440; // @[control.scala 438:19 296:35]
  wire  _GEN_1482 = 6'h9 == state ? ofm_recv_task_enable : _GEN_1441; // @[control.scala 438:19 358:39]
  wire  _GEN_1483 = 6'h9 == state ? first_ofm_recv_stop : _GEN_1442; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1484 = 6'h9 == state ? ofm_addr_fmbase : _GEN_1443; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1485 = 6'h9 == state ? ofm_addr_offset : _GEN_1444; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1486 = 6'h9 == state ? ofm_recv_len : _GEN_1445; // @[control.scala 438:19 367:31]
  wire  _GEN_1487 = 6'h9 == state ? wgt_send_task_enable : _GEN_1446; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1488 = 6'h9 == state ? wgt_addr_send : _GEN_1447; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1489 = 6'h9 == state ? wgt_addr_read : _GEN_1448; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1490 = 6'h9 == state ? iter_ifm_post : _GEN_1449; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1491 = 6'h9 == state ? iter_div_post : _GEN_1450; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1492 = 6'h9 == state ? iter_ofm_post : _GEN_1451; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1493 = 6'h9 == state ? iter_ifm_pre : _GEN_1452; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1494 = 6'h9 == state ? iter_div_pre : _GEN_1453; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1495 = 6'h9 == state ? iter_ofm_pre : _GEN_1454; // @[control.scala 438:19 194:31]
  wire  _GEN_1496 = 6'h9 == state ? ifm_send_task_enable : _GEN_1455; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1497 = 6'h9 == state ? ifm_addr_fmbase : _GEN_1456; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1498 = 6'h9 == state ? ifm_addr_offset : _GEN_1457; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1499 = 6'h9 == state ? ifm_send_len : _GEN_1458; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1500 = 6'h9 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1459; // @[control.scala 438:19 425:46]
  wire [25:0] _GEN_1501 = 6'h9 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1460; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1502 = 6'h9 == state ? weight_sel : _GEN_1461; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1503 = 6'h9 == state ? bia_addr_read : _GEN_1462; // @[control.scala 438:19 181:32]
  wire  _GEN_1504 = 6'h9 == state ? wgt_ddr_read_en : _GEN_1463; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1505 = 6'h9 == state ? reg_t_6 : _GEN_1464; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1506 = 6'h9 == state ? reg_t_7 : _GEN_1465; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1507 = 6'h9 == state ? pool_cnt : _GEN_1466; // @[control.scala 438:19 290:27]
  wire  _GEN_1508 = 6'h9 == state ? ifm_sel : _GEN_1467; // @[control.scala 438:19 379:24]
  wire  _GEN_1509 = 6'h9 == state ? resize_load_t : _GEN_1468; // @[control.scala 438:19 420:32]
  wire  _GEN_1510 = 6'h9 == state ? yolo_finish : _GEN_1469; // @[control.scala 438:19 40:28]
  wire  _GEN_1511 = 6'h9 == state ? conv_finish : _GEN_1470; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1512 = 6'h8 == state ? _ifm_addr_fmbase_T : _GEN_1497; // @[control.scala 438:19 540:29]
  wire [31:0] _GEN_1513 = 6'h8 == state ? _GEN_45 : _GEN_1498; // @[control.scala 438:19]
  wire [31:0] _GEN_1514 = 6'h8 == state ? _GEN_46 : _GEN_1499; // @[control.scala 438:19]
  wire [9:0] _GEN_1515 = 6'h8 == state ? _GEN_47 : _GEN_1500; // @[control.scala 438:19]
  wire [31:0] _GEN_1516 = 6'h8 == state ? _GEN_48 : _GEN_1471; // @[control.scala 438:19]
  wire [5:0] _GEN_1517 = 6'h8 == state ? 6'h9 : _GEN_1472; // @[control.scala 438:19 600:19]
  wire  _GEN_1518 = 6'h8 == state ? last_buf_sel : _GEN_1473; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1519 = 6'h8 == state ? reg_task : _GEN_1474; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1520 = 6'h8 == state ? reg_t_4 : _GEN_1475; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1521 = 6'h8 == state ? reg_t_5 : _GEN_1476; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1522 = 6'h8 == state ? reg_t_3 : _GEN_1477; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1523 = 6'h8 == state ? reg_t_0 : _GEN_1478; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1524 = 6'h8 == state ? cnt_t : _GEN_1479; // @[control.scala 438:19 163:24]
  wire  _GEN_1525 = 6'h8 == state ? bottleneck_transfer : _GEN_1480; // @[control.scala 438:19 295:38]
  wire  _GEN_1526 = 6'h8 == state ? bottleneck_ready : _GEN_1481; // @[control.scala 438:19 296:35]
  wire  _GEN_1527 = 6'h8 == state ? ofm_recv_task_enable : _GEN_1482; // @[control.scala 438:19 358:39]
  wire  _GEN_1528 = 6'h8 == state ? first_ofm_recv_stop : _GEN_1483; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1529 = 6'h8 == state ? ofm_addr_fmbase : _GEN_1484; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1530 = 6'h8 == state ? ofm_addr_offset : _GEN_1485; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1531 = 6'h8 == state ? ofm_recv_len : _GEN_1486; // @[control.scala 438:19 367:31]
  wire  _GEN_1532 = 6'h8 == state ? wgt_send_task_enable : _GEN_1487; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1533 = 6'h8 == state ? wgt_addr_send : _GEN_1488; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1534 = 6'h8 == state ? wgt_addr_read : _GEN_1489; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1535 = 6'h8 == state ? iter_ifm_post : _GEN_1490; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1536 = 6'h8 == state ? iter_div_post : _GEN_1491; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1537 = 6'h8 == state ? iter_ofm_post : _GEN_1492; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1538 = 6'h8 == state ? iter_ifm_pre : _GEN_1493; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1539 = 6'h8 == state ? iter_div_pre : _GEN_1494; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1540 = 6'h8 == state ? iter_ofm_pre : _GEN_1495; // @[control.scala 438:19 194:31]
  wire  _GEN_1541 = 6'h8 == state ? ifm_send_task_enable : _GEN_1496; // @[control.scala 438:19 357:39]
  wire [25:0] _GEN_1542 = 6'h8 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1501; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1543 = 6'h8 == state ? weight_sel : _GEN_1502; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1544 = 6'h8 == state ? bia_addr_read : _GEN_1503; // @[control.scala 438:19 181:32]
  wire  _GEN_1545 = 6'h8 == state ? wgt_ddr_read_en : _GEN_1504; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1546 = 6'h8 == state ? reg_t_6 : _GEN_1505; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1547 = 6'h8 == state ? reg_t_7 : _GEN_1506; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1548 = 6'h8 == state ? pool_cnt : _GEN_1507; // @[control.scala 438:19 290:27]
  wire  _GEN_1549 = 6'h8 == state ? ifm_sel : _GEN_1508; // @[control.scala 438:19 379:24]
  wire  _GEN_1550 = 6'h8 == state ? resize_load_t : _GEN_1509; // @[control.scala 438:19 420:32]
  wire  _GEN_1551 = 6'h8 == state ? yolo_finish : _GEN_1510; // @[control.scala 438:19 40:28]
  wire  _GEN_1552 = 6'h8 == state ? conv_finish : _GEN_1511; // @[control.scala 438:19 71:30]
  wire  _GEN_1553 = 6'h7 == state ? _T_13 : _GEN_1541; // @[control.scala 438:19]
  wire [5:0] _GEN_1554 = 6'h7 == state ? {{2'd0}, _GEN_18} : _GEN_1517; // @[control.scala 438:19]
  wire [31:0] _GEN_1555 = 6'h7 == state ? ifm_addr_fmbase : _GEN_1512; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1556 = 6'h7 == state ? ifm_addr_offset : _GEN_1513; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1557 = 6'h7 == state ? ifm_send_len : _GEN_1514; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1558 = 6'h7 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1515; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1559 = 6'h7 == state ? reg_static : _GEN_1516; // @[control.scala 438:19 161:29]
  wire  _GEN_1560 = 6'h7 == state ? last_buf_sel : _GEN_1518; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1561 = 6'h7 == state ? reg_task : _GEN_1519; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1562 = 6'h7 == state ? reg_t_4 : _GEN_1520; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1563 = 6'h7 == state ? reg_t_5 : _GEN_1521; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1564 = 6'h7 == state ? reg_t_3 : _GEN_1522; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1565 = 6'h7 == state ? reg_t_0 : _GEN_1523; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1566 = 6'h7 == state ? cnt_t : _GEN_1524; // @[control.scala 438:19 163:24]
  wire  _GEN_1567 = 6'h7 == state ? bottleneck_transfer : _GEN_1525; // @[control.scala 438:19 295:38]
  wire  _GEN_1568 = 6'h7 == state ? bottleneck_ready : _GEN_1526; // @[control.scala 438:19 296:35]
  wire  _GEN_1569 = 6'h7 == state ? ofm_recv_task_enable : _GEN_1527; // @[control.scala 438:19 358:39]
  wire  _GEN_1570 = 6'h7 == state ? first_ofm_recv_stop : _GEN_1528; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1571 = 6'h7 == state ? ofm_addr_fmbase : _GEN_1529; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1572 = 6'h7 == state ? ofm_addr_offset : _GEN_1530; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1573 = 6'h7 == state ? ofm_recv_len : _GEN_1531; // @[control.scala 438:19 367:31]
  wire  _GEN_1574 = 6'h7 == state ? wgt_send_task_enable : _GEN_1532; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1575 = 6'h7 == state ? wgt_addr_send : _GEN_1533; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1576 = 6'h7 == state ? wgt_addr_read : _GEN_1534; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1577 = 6'h7 == state ? iter_ifm_post : _GEN_1535; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1578 = 6'h7 == state ? iter_div_post : _GEN_1536; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1579 = 6'h7 == state ? iter_ofm_post : _GEN_1537; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1580 = 6'h7 == state ? iter_ifm_pre : _GEN_1538; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1581 = 6'h7 == state ? iter_div_pre : _GEN_1539; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1582 = 6'h7 == state ? iter_ofm_pre : _GEN_1540; // @[control.scala 438:19 194:31]
  wire [25:0] _GEN_1583 = 6'h7 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1542; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1584 = 6'h7 == state ? weight_sel : _GEN_1543; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1585 = 6'h7 == state ? bia_addr_read : _GEN_1544; // @[control.scala 438:19 181:32]
  wire  _GEN_1586 = 6'h7 == state ? wgt_ddr_read_en : _GEN_1545; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1587 = 6'h7 == state ? reg_t_6 : _GEN_1546; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1588 = 6'h7 == state ? reg_t_7 : _GEN_1547; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1589 = 6'h7 == state ? pool_cnt : _GEN_1548; // @[control.scala 438:19 290:27]
  wire  _GEN_1590 = 6'h7 == state ? ifm_sel : _GEN_1549; // @[control.scala 438:19 379:24]
  wire  _GEN_1591 = 6'h7 == state ? resize_load_t : _GEN_1550; // @[control.scala 438:19 420:32]
  wire  _GEN_1592 = 6'h7 == state ? yolo_finish : _GEN_1551; // @[control.scala 438:19 40:28]
  wire  _GEN_1593 = 6'h7 == state ? conv_finish : _GEN_1552; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_1594 = 6'h6 == state ? {{3'd0}, _GEN_16} : _GEN_1554; // @[control.scala 438:19]
  wire  _GEN_1595 = 6'h6 == state ? ifm_send_task_enable : _GEN_1553; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1596 = 6'h6 == state ? ifm_addr_fmbase : _GEN_1555; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1597 = 6'h6 == state ? ifm_addr_offset : _GEN_1556; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1598 = 6'h6 == state ? ifm_send_len : _GEN_1557; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1599 = 6'h6 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1558; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1600 = 6'h6 == state ? reg_static : _GEN_1559; // @[control.scala 438:19 161:29]
  wire  _GEN_1601 = 6'h6 == state ? last_buf_sel : _GEN_1560; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1602 = 6'h6 == state ? reg_task : _GEN_1561; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1603 = 6'h6 == state ? reg_t_4 : _GEN_1562; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1604 = 6'h6 == state ? reg_t_5 : _GEN_1563; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1605 = 6'h6 == state ? reg_t_3 : _GEN_1564; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1606 = 6'h6 == state ? reg_t_0 : _GEN_1565; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1607 = 6'h6 == state ? cnt_t : _GEN_1566; // @[control.scala 438:19 163:24]
  wire  _GEN_1608 = 6'h6 == state ? bottleneck_transfer : _GEN_1567; // @[control.scala 438:19 295:38]
  wire  _GEN_1609 = 6'h6 == state ? bottleneck_ready : _GEN_1568; // @[control.scala 438:19 296:35]
  wire  _GEN_1610 = 6'h6 == state ? ofm_recv_task_enable : _GEN_1569; // @[control.scala 438:19 358:39]
  wire  _GEN_1611 = 6'h6 == state ? first_ofm_recv_stop : _GEN_1570; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1612 = 6'h6 == state ? ofm_addr_fmbase : _GEN_1571; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1613 = 6'h6 == state ? ofm_addr_offset : _GEN_1572; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1614 = 6'h6 == state ? ofm_recv_len : _GEN_1573; // @[control.scala 438:19 367:31]
  wire  _GEN_1615 = 6'h6 == state ? wgt_send_task_enable : _GEN_1574; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1616 = 6'h6 == state ? wgt_addr_send : _GEN_1575; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1617 = 6'h6 == state ? wgt_addr_read : _GEN_1576; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1618 = 6'h6 == state ? iter_ifm_post : _GEN_1577; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1619 = 6'h6 == state ? iter_div_post : _GEN_1578; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1620 = 6'h6 == state ? iter_ofm_post : _GEN_1579; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1621 = 6'h6 == state ? iter_ifm_pre : _GEN_1580; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1622 = 6'h6 == state ? iter_div_pre : _GEN_1581; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1623 = 6'h6 == state ? iter_ofm_pre : _GEN_1582; // @[control.scala 438:19 194:31]
  wire [25:0] _GEN_1624 = 6'h6 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1583; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1625 = 6'h6 == state ? weight_sel : _GEN_1584; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1626 = 6'h6 == state ? bia_addr_read : _GEN_1585; // @[control.scala 438:19 181:32]
  wire  _GEN_1627 = 6'h6 == state ? wgt_ddr_read_en : _GEN_1586; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1628 = 6'h6 == state ? reg_t_6 : _GEN_1587; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1629 = 6'h6 == state ? reg_t_7 : _GEN_1588; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1630 = 6'h6 == state ? pool_cnt : _GEN_1589; // @[control.scala 438:19 290:27]
  wire  _GEN_1631 = 6'h6 == state ? ifm_sel : _GEN_1590; // @[control.scala 438:19 379:24]
  wire  _GEN_1632 = 6'h6 == state ? resize_load_t : _GEN_1591; // @[control.scala 438:19 420:32]
  wire  _GEN_1633 = 6'h6 == state ? yolo_finish : _GEN_1592; // @[control.scala 438:19 40:28]
  wire  _GEN_1634 = 6'h6 == state ? conv_finish : _GEN_1593; // @[control.scala 438:19 71:30]
  wire [4:0] _GEN_1635 = 6'h5 == state ? _GEN_2 : _GEN_1607; // @[control.scala 438:19]
  wire [5:0] _GEN_1636 = 6'h5 == state ? _GEN_10 : _GEN_1594; // @[control.scala 438:19]
  wire [31:0] _GEN_1637 = 6'h5 == state ? _GEN_11 : _GEN_1606; // @[control.scala 438:19]
  wire [31:0] _GEN_1638 = 6'h5 == state ? _GEN_12 : reg_t_1; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1639 = 6'h5 == state ? _GEN_13 : reg_t_2; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1640 = 6'h5 == state ? _GEN_14 : reg_t_9; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1641 = 6'h5 == state ? _GEN_15 : reg_t_10; // @[control.scala 438:19 160:37]
  wire  _GEN_1642 = 6'h5 == state ? ifm_send_task_enable : _GEN_1595; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1643 = 6'h5 == state ? ifm_addr_fmbase : _GEN_1596; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1644 = 6'h5 == state ? ifm_addr_offset : _GEN_1597; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1645 = 6'h5 == state ? ifm_send_len : _GEN_1598; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1646 = 6'h5 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1599; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1647 = 6'h5 == state ? reg_static : _GEN_1600; // @[control.scala 438:19 161:29]
  wire  _GEN_1648 = 6'h5 == state ? last_buf_sel : _GEN_1601; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1649 = 6'h5 == state ? reg_task : _GEN_1602; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1650 = 6'h5 == state ? reg_t_4 : _GEN_1603; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1651 = 6'h5 == state ? reg_t_5 : _GEN_1604; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1652 = 6'h5 == state ? reg_t_3 : _GEN_1605; // @[control.scala 438:19 160:37]
  wire  _GEN_1653 = 6'h5 == state ? bottleneck_transfer : _GEN_1608; // @[control.scala 438:19 295:38]
  wire  _GEN_1654 = 6'h5 == state ? bottleneck_ready : _GEN_1609; // @[control.scala 438:19 296:35]
  wire  _GEN_1655 = 6'h5 == state ? ofm_recv_task_enable : _GEN_1610; // @[control.scala 438:19 358:39]
  wire  _GEN_1656 = 6'h5 == state ? first_ofm_recv_stop : _GEN_1611; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1657 = 6'h5 == state ? ofm_addr_fmbase : _GEN_1612; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1658 = 6'h5 == state ? ofm_addr_offset : _GEN_1613; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1659 = 6'h5 == state ? ofm_recv_len : _GEN_1614; // @[control.scala 438:19 367:31]
  wire  _GEN_1660 = 6'h5 == state ? wgt_send_task_enable : _GEN_1615; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1661 = 6'h5 == state ? wgt_addr_send : _GEN_1616; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1662 = 6'h5 == state ? wgt_addr_read : _GEN_1617; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1663 = 6'h5 == state ? iter_ifm_post : _GEN_1618; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1664 = 6'h5 == state ? iter_div_post : _GEN_1619; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1665 = 6'h5 == state ? iter_ofm_post : _GEN_1620; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1666 = 6'h5 == state ? iter_ifm_pre : _GEN_1621; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1667 = 6'h5 == state ? iter_div_pre : _GEN_1622; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1668 = 6'h5 == state ? iter_ofm_pre : _GEN_1623; // @[control.scala 438:19 194:31]
  wire [25:0] _GEN_1669 = 6'h5 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1624; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1670 = 6'h5 == state ? weight_sel : _GEN_1625; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1671 = 6'h5 == state ? bia_addr_read : _GEN_1626; // @[control.scala 438:19 181:32]
  wire  _GEN_1672 = 6'h5 == state ? wgt_ddr_read_en : _GEN_1627; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1673 = 6'h5 == state ? reg_t_6 : _GEN_1628; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1674 = 6'h5 == state ? reg_t_7 : _GEN_1629; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1675 = 6'h5 == state ? pool_cnt : _GEN_1630; // @[control.scala 438:19 290:27]
  wire  _GEN_1676 = 6'h5 == state ? ifm_sel : _GEN_1631; // @[control.scala 438:19 379:24]
  wire  _GEN_1677 = 6'h5 == state ? resize_load_t : _GEN_1632; // @[control.scala 438:19 420:32]
  wire  _GEN_1678 = 6'h5 == state ? yolo_finish : _GEN_1633; // @[control.scala 438:19 40:28]
  wire  _GEN_1679 = 6'h5 == state ? conv_finish : _GEN_1634; // @[control.scala 438:19 71:30]
  wire [31:0] _GEN_1680 = 6'h4 == state ? wgt_ddr_base_addr : _GEN_1650; // @[control.scala 438:19 498:22]
  wire [31:0] _GEN_1681 = 6'h4 == state ? {{12'd0}, _reg_t_5_T_6} : _GEN_1651; // @[control.scala 438:19 499:22]
  wire [31:0] _GEN_1682 = 6'h4 == state ? 32'h205 : _GEN_1637; // @[control.scala 438:19 500:22]
  wire [4:0] _GEN_1683 = 6'h4 == state ? 5'h0 : _GEN_1635; // @[control.scala 438:19 501:19]
  wire [5:0] _GEN_1684 = 6'h4 == state ? 6'h5 : _GEN_1636; // @[control.scala 438:19 502:19]
  wire [31:0] _GEN_1685 = 6'h4 == state ? reg_t_1 : _GEN_1638; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1686 = 6'h4 == state ? reg_t_2 : _GEN_1639; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1687 = 6'h4 == state ? reg_t_9 : _GEN_1640; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1688 = 6'h4 == state ? reg_t_10 : _GEN_1641; // @[control.scala 438:19 160:37]
  wire  _GEN_1689 = 6'h4 == state ? ifm_send_task_enable : _GEN_1642; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1690 = 6'h4 == state ? ifm_addr_fmbase : _GEN_1643; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1691 = 6'h4 == state ? ifm_addr_offset : _GEN_1644; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1692 = 6'h4 == state ? ifm_send_len : _GEN_1645; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1693 = 6'h4 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1646; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1694 = 6'h4 == state ? reg_static : _GEN_1647; // @[control.scala 438:19 161:29]
  wire  _GEN_1695 = 6'h4 == state ? last_buf_sel : _GEN_1648; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1696 = 6'h4 == state ? reg_task : _GEN_1649; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1697 = 6'h4 == state ? reg_t_3 : _GEN_1652; // @[control.scala 438:19 160:37]
  wire  _GEN_1698 = 6'h4 == state ? bottleneck_transfer : _GEN_1653; // @[control.scala 438:19 295:38]
  wire  _GEN_1699 = 6'h4 == state ? bottleneck_ready : _GEN_1654; // @[control.scala 438:19 296:35]
  wire  _GEN_1700 = 6'h4 == state ? ofm_recv_task_enable : _GEN_1655; // @[control.scala 438:19 358:39]
  wire  _GEN_1701 = 6'h4 == state ? first_ofm_recv_stop : _GEN_1656; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1702 = 6'h4 == state ? ofm_addr_fmbase : _GEN_1657; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1703 = 6'h4 == state ? ofm_addr_offset : _GEN_1658; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1704 = 6'h4 == state ? ofm_recv_len : _GEN_1659; // @[control.scala 438:19 367:31]
  wire  _GEN_1705 = 6'h4 == state ? wgt_send_task_enable : _GEN_1660; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1706 = 6'h4 == state ? wgt_addr_send : _GEN_1661; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1707 = 6'h4 == state ? wgt_addr_read : _GEN_1662; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1708 = 6'h4 == state ? iter_ifm_post : _GEN_1663; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1709 = 6'h4 == state ? iter_div_post : _GEN_1664; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1710 = 6'h4 == state ? iter_ofm_post : _GEN_1665; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1711 = 6'h4 == state ? iter_ifm_pre : _GEN_1666; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1712 = 6'h4 == state ? iter_div_pre : _GEN_1667; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1713 = 6'h4 == state ? iter_ofm_pre : _GEN_1668; // @[control.scala 438:19 194:31]
  wire [25:0] _GEN_1714 = 6'h4 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1669; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1715 = 6'h4 == state ? weight_sel : _GEN_1670; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1716 = 6'h4 == state ? bia_addr_read : _GEN_1671; // @[control.scala 438:19 181:32]
  wire  _GEN_1717 = 6'h4 == state ? wgt_ddr_read_en : _GEN_1672; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1718 = 6'h4 == state ? reg_t_6 : _GEN_1673; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1719 = 6'h4 == state ? reg_t_7 : _GEN_1674; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1720 = 6'h4 == state ? pool_cnt : _GEN_1675; // @[control.scala 438:19 290:27]
  wire  _GEN_1721 = 6'h4 == state ? ifm_sel : _GEN_1676; // @[control.scala 438:19 379:24]
  wire  _GEN_1722 = 6'h4 == state ? resize_load_t : _GEN_1677; // @[control.scala 438:19 420:32]
  wire  _GEN_1723 = 6'h4 == state ? yolo_finish : _GEN_1678; // @[control.scala 438:19 40:28]
  wire  _GEN_1724 = 6'h4 == state ? conv_finish : _GEN_1679; // @[control.scala 438:19 71:30]
  wire [5:0] _GEN_1725 = 6'h3 == state ? {{3'd0}, _GEN_8} : _GEN_1684; // @[control.scala 438:19]
  wire [31:0] _GEN_1726 = 6'h3 == state ? reg_t_4 : _GEN_1680; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1727 = 6'h3 == state ? reg_t_5 : _GEN_1681; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1728 = 6'h3 == state ? reg_t_0 : _GEN_1682; // @[control.scala 438:19 160:37]
  wire [4:0] _GEN_1729 = 6'h3 == state ? cnt_t : _GEN_1683; // @[control.scala 438:19 163:24]
  wire [31:0] _GEN_1730 = 6'h3 == state ? reg_t_1 : _GEN_1685; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1731 = 6'h3 == state ? reg_t_2 : _GEN_1686; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1732 = 6'h3 == state ? reg_t_9 : _GEN_1687; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1733 = 6'h3 == state ? reg_t_10 : _GEN_1688; // @[control.scala 438:19 160:37]
  wire  _GEN_1734 = 6'h3 == state ? ifm_send_task_enable : _GEN_1689; // @[control.scala 438:19 357:39]
  wire [31:0] _GEN_1735 = 6'h3 == state ? ifm_addr_fmbase : _GEN_1690; // @[control.scala 438:19 362:34]
  wire [31:0] _GEN_1736 = 6'h3 == state ? ifm_addr_offset : _GEN_1691; // @[control.scala 438:19 363:34]
  wire [31:0] _GEN_1737 = 6'h3 == state ? ifm_send_len : _GEN_1692; // @[control.scala 438:19 364:31]
  wire [9:0] _GEN_1738 = 6'h3 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1693; // @[control.scala 438:19 425:46]
  wire [31:0] _GEN_1739 = 6'h3 == state ? reg_static : _GEN_1694; // @[control.scala 438:19 161:29]
  wire  _GEN_1740 = 6'h3 == state ? last_buf_sel : _GEN_1695; // @[control.scala 438:19 182:31]
  wire [31:0] _GEN_1741 = 6'h3 == state ? reg_task : _GEN_1696; // @[control.scala 438:19 162:27]
  wire [31:0] _GEN_1742 = 6'h3 == state ? reg_t_3 : _GEN_1697; // @[control.scala 438:19 160:37]
  wire  _GEN_1743 = 6'h3 == state ? bottleneck_transfer : _GEN_1698; // @[control.scala 438:19 295:38]
  wire  _GEN_1744 = 6'h3 == state ? bottleneck_ready : _GEN_1699; // @[control.scala 438:19 296:35]
  wire  _GEN_1745 = 6'h3 == state ? ofm_recv_task_enable : _GEN_1700; // @[control.scala 438:19 358:39]
  wire  _GEN_1746 = 6'h3 == state ? first_ofm_recv_stop : _GEN_1701; // @[control.scala 438:19 422:38]
  wire [31:0] _GEN_1747 = 6'h3 == state ? ofm_addr_fmbase : _GEN_1702; // @[control.scala 438:19 365:34]
  wire [31:0] _GEN_1748 = 6'h3 == state ? ofm_addr_offset : _GEN_1703; // @[control.scala 438:19 366:34]
  wire [31:0] _GEN_1749 = 6'h3 == state ? ofm_recv_len : _GEN_1704; // @[control.scala 438:19 367:31]
  wire  _GEN_1750 = 6'h3 == state ? wgt_send_task_enable : _GEN_1705; // @[control.scala 438:19 359:39]
  wire [31:0] _GEN_1751 = 6'h3 == state ? wgt_addr_send : _GEN_1706; // @[control.scala 438:19 178:32]
  wire [15:0] _GEN_1752 = 6'h3 == state ? wgt_addr_read : _GEN_1707; // @[control.scala 438:19 179:32]
  wire [12:0] _GEN_1753 = 6'h3 == state ? iter_ifm_post : _GEN_1708; // @[control.scala 438:19 196:32]
  wire [12:0] _GEN_1754 = 6'h3 == state ? iter_div_post : _GEN_1709; // @[control.scala 438:19 198:32]
  wire [12:0] _GEN_1755 = 6'h3 == state ? iter_ofm_post : _GEN_1710; // @[control.scala 438:19 197:32]
  wire [12:0] _GEN_1756 = 6'h3 == state ? iter_ifm_pre : _GEN_1711; // @[control.scala 438:19 192:31]
  wire [12:0] _GEN_1757 = 6'h3 == state ? iter_div_pre : _GEN_1712; // @[control.scala 438:19 195:31]
  wire [12:0] _GEN_1758 = 6'h3 == state ? iter_ofm_pre : _GEN_1713; // @[control.scala 438:19 194:31]
  wire [25:0] _GEN_1759 = 6'h3 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1714; // @[control.scala 438:19 180:34]
  wire [2:0] _GEN_1760 = 6'h3 == state ? weight_sel : _GEN_1715; // @[control.scala 438:19 274:27]
  wire [15:0] _GEN_1761 = 6'h3 == state ? bia_addr_read : _GEN_1716; // @[control.scala 438:19 181:32]
  wire  _GEN_1762 = 6'h3 == state ? wgt_ddr_read_en : _GEN_1717; // @[control.scala 438:19 424:32]
  wire [31:0] _GEN_1763 = 6'h3 == state ? reg_t_6 : _GEN_1718; // @[control.scala 438:19 160:37]
  wire [31:0] _GEN_1764 = 6'h3 == state ? reg_t_7 : _GEN_1719; // @[control.scala 438:19 160:37]
  wire [1:0] _GEN_1765 = 6'h3 == state ? pool_cnt : _GEN_1720; // @[control.scala 438:19 290:27]
  wire  _GEN_1766 = 6'h3 == state ? ifm_sel : _GEN_1721; // @[control.scala 438:19 379:24]
  wire  _GEN_1767 = 6'h3 == state ? resize_load_t : _GEN_1722; // @[control.scala 438:19 420:32]
  wire  _GEN_1768 = 6'h3 == state ? yolo_finish : _GEN_1723; // @[control.scala 438:19 40:28]
  wire  _GEN_1769 = 6'h3 == state ? conv_finish : _GEN_1724; // @[control.scala 438:19 71:30]
  wire [9:0] _GEN_1783 = 6'h2 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1738; // @[control.scala 438:19 425:46]
  wire [25:0] _GEN_1804 = 6'h2 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1759; // @[control.scala 438:19 180:34]
  wire [9:0] _GEN_1842 = 6'h1 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1783; // @[control.scala 438:19 425:46]
  wire [25:0] _GEN_1852 = 6'h1 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1804; // @[control.scala 438:19 180:34]
  wire [9:0] _GEN_1890 = 6'h0 == state ? {{2'd0}, the_number_of_row_transferred} : _GEN_1842; // @[control.scala 438:19 425:46]
  wire [25:0] _GEN_1899 = 6'h0 == state ? {{10'd0}, wgt_addr_read_t} : _GEN_1852; // @[control.scala 438:19 180:34]
  wire [2:0] _conv_in_c2f_T_2 = _c2f_shortcut_T_1 ? 3'h6 : 3'h3; // @[Mux.scala 101:16]
  wire [2:0] _conv_in_c2f_T_3 = _c2f_shortcut_T ? 3'h6 : _conv_in_c2f_T_2; // @[Mux.scala 101:16]
  wire [1:0] conv_in_c2f = _conv_in_c2f_T_3[1:0]; // @[control.scala 1299:27 1300:17]
  wire [2:0] _cur_conv_in_c2f_T = {conv_in_c2f, 1'h0}; // @[control.scala 1301:46]
  wire [2:0] cur_conv_in_c2f = 3'h2 + _cur_conv_in_c2f_T; // @[control.scala 1301:31]
  wire [2:0] _everu_layer_conv_number_T_3 = 3'h1 == current_model_code ? cur_conv_in_c2f : {{2'd0}, 3'h0 ==
    current_model_code}; // @[Mux.scala 81:58]
  wire [2:0] _everu_layer_conv_number_T_5 = 3'h2 == current_model_code ? 3'h2 : _everu_layer_conv_number_T_3; // @[Mux.scala 81:58]
  wire [2:0] _everu_layer_conv_number_T_7 = 3'h3 == current_model_code ? 3'h3 : _everu_layer_conv_number_T_5; // @[Mux.scala 81:58]
  wire [2:0] _everu_layer_conv_number_T_9 = 3'h4 == current_model_code ? 3'h3 : _everu_layer_conv_number_T_7; // @[Mux.scala 81:58]
  reg  conv_cnt; // @[control.scala 1305:25]
  reg [6:0] base; // @[control.scala 1309:21]
  reg [6:0] cnt_layer; // @[control.scala 1312:28]
  wire [4:0] everu_layer_conv_number = {{2'd0}, _everu_layer_conv_number_T_9}; // @[control.scala 1302:39 1303:29]
  wire [6:0] _GEN_2858 = {{2'd0}, everu_layer_conv_number}; // @[control.scala 1313:83]
  wire [6:0] _base_T_2 = base + _GEN_2858; // @[control.scala 1313:83]
  wire [6:0] _GEN_2859 = {{6'd0}, conv_cnt}; // @[control.scala 1314:20]
  wire [6:0] _cnt_layer_T_1 = base + _GEN_2859; // @[control.scala 1314:20]
  wire [15:0] _GEN_1905 = 7'h66 == cnt_layer ? 16'h4868 : conv_scale; // @[control.scala 1315:23 2475:25 112:28]
  wire [3:0] _GEN_1906 = 7'h66 == cnt_layer ? 4'h7 : conv_shift; // @[control.scala 1315:23 2476:25 113:29]
  wire [7:0] _GEN_1907 = 7'h66 == cnt_layer ? 8'h0 : zp_in; // @[control.scala 1315:23 114:24 2477:25]
  wire [7:0] _GEN_1908 = 7'h66 == cnt_layer ? 8'h79 : zp_out; // @[control.scala 1315:23 115:25 2478:25]
  wire [31:0] _GEN_1909 = 7'h66 == cnt_layer ? 32'h3f05b3e5 : scale_B_act; // @[control.scala 1315:23 2479:25 117:30]
  wire [31:0] _GEN_1910 = 7'h66 == cnt_layer ? 32'h42122c8f : scale_A_act; // @[control.scala 1315:23 2480:25 118:30]
  wire [7:0] _GEN_1911 = 7'h66 == cnt_layer ? 8'ha : zp_act; // @[control.scala 1315:23 116:25 2481:25]
  wire [31:0] _GEN_1912 = 7'h66 == cnt_layer ? 32'h22cb0000 : wgt_ddr_base_addr; // @[control.scala 1315:23 2482:31 369:36]
  wire [31:0] _GEN_1913 = 7'h66 == cnt_layer ? 32'h22d2b000 : bia_ddr_base_addr; // @[control.scala 1315:23 2483:31 370:36]
  wire [15:0] _GEN_1914 = 7'h65 == cnt_layer ? 16'h5a61 : _GEN_1905; // @[control.scala 1315:23 2464:25]
  wire [3:0] _GEN_1915 = 7'h65 == cnt_layer ? 4'h7 : _GEN_1906; // @[control.scala 1315:23 2465:25]
  wire [7:0] _GEN_1916 = 7'h65 == cnt_layer ? 8'h3 : _GEN_1907; // @[control.scala 1315:23 2466:25]
  wire [7:0] _GEN_1917 = 7'h65 == cnt_layer ? 8'h3b : _GEN_1908; // @[control.scala 1315:23 2467:25]
  wire [31:0] _GEN_1918 = 7'h65 == cnt_layer ? 32'h3fbe3417 : _GEN_1909; // @[control.scala 1315:23 2468:25]
  wire [31:0] _GEN_1919 = 7'h65 == cnt_layer ? 32'h3fa16942 : _GEN_1910; // @[control.scala 1315:23 2469:25]
  wire [7:0] _GEN_1920 = 7'h65 == cnt_layer ? 8'h0 : _GEN_1911; // @[control.scala 1315:23 2470:25]
  wire [31:0] _GEN_1921 = 7'h65 == cnt_layer ? 32'h22c68000 : _GEN_1912; // @[control.scala 1315:23 2471:31]
  wire [31:0] _GEN_1922 = 7'h65 == cnt_layer ? 32'h22d2a800 : _GEN_1913; // @[control.scala 1315:23 2472:31]
  wire [15:0] _GEN_1923 = 7'h64 == cnt_layer ? 16'h4672 : _GEN_1914; // @[control.scala 1315:23 2453:25]
  wire [3:0] _GEN_1924 = 7'h64 == cnt_layer ? 4'h7 : _GEN_1915; // @[control.scala 1315:23 2454:25]
  wire [7:0] _GEN_1925 = 7'h64 == cnt_layer ? 8'h3 : _GEN_1916; // @[control.scala 1315:23 2455:25]
  wire [7:0] _GEN_1926 = 7'h64 == cnt_layer ? 8'h5e : _GEN_1917; // @[control.scala 1315:23 2456:25]
  wire [31:0] _GEN_1927 = 7'h64 == cnt_layer ? 32'h3ec30b3e : _GEN_1918; // @[control.scala 1315:23 2457:25]
  wire [31:0] _GEN_1928 = 7'h64 == cnt_layer ? 32'h411c604b : _GEN_1919; // @[control.scala 1315:23 2458:25]
  wire [7:0] _GEN_1929 = 7'h64 == cnt_layer ? 8'h3 : _GEN_1920; // @[control.scala 1315:23 2459:25]
  wire [31:0] _GEN_1930 = 7'h64 == cnt_layer ? 32'h22c20000 : _GEN_1921; // @[control.scala 1315:23 2460:31]
  wire [31:0] _GEN_1931 = 7'h64 == cnt_layer ? 32'h22d2a000 : _GEN_1922; // @[control.scala 1315:23 2461:31]
  wire [15:0] _GEN_1932 = 7'h63 == cnt_layer ? 16'h5aa9 : _GEN_1923; // @[control.scala 1315:23 2441:25]
  wire [3:0] _GEN_1933 = 7'h63 == cnt_layer ? 4'h7 : _GEN_1924; // @[control.scala 1315:23 2442:25]
  wire [7:0] _GEN_1934 = 7'h63 == cnt_layer ? 8'h0 : _GEN_1925; // @[control.scala 1315:23 2443:25]
  wire [7:0] _GEN_1935 = 7'h63 == cnt_layer ? 8'h79 : _GEN_1926; // @[control.scala 1315:23 2444:25]
  wire [31:0] _GEN_1936 = 7'h63 == cnt_layer ? 32'h3eff5cc1 : _GEN_1927; // @[control.scala 1315:23 2445:25]
  wire [31:0] _GEN_1937 = 7'h63 == cnt_layer ? 32'h4220d9d7 : _GEN_1928; // @[control.scala 1315:23 2446:25]
  wire [7:0] _GEN_1938 = 7'h63 == cnt_layer ? 8'hb : _GEN_1929; // @[control.scala 1315:23 2447:25]
  wire [31:0] _GEN_1939 = 7'h63 == cnt_layer ? 32'h22bd8000 : _GEN_1930; // @[control.scala 1315:23 2448:31]
  wire [31:0] _GEN_1940 = 7'h63 == cnt_layer ? 32'h22d29800 : _GEN_1931; // @[control.scala 1315:23 2449:31]
  wire [15:0] _GEN_1941 = 7'h62 == cnt_layer ? 16'h4c1a : _GEN_1932; // @[control.scala 1315:23 2430:25]
  wire [3:0] _GEN_1942 = 7'h62 == cnt_layer ? 4'h7 : _GEN_1933; // @[control.scala 1315:23 2431:25]
  wire [7:0] _GEN_1943 = 7'h62 == cnt_layer ? 8'h3 : _GEN_1934; // @[control.scala 1315:23 2432:25]
  wire [7:0] _GEN_1944 = 7'h62 == cnt_layer ? 8'h3d : _GEN_1935; // @[control.scala 1315:23 2433:25]
  wire [31:0] _GEN_1945 = 7'h62 == cnt_layer ? 32'h4014cdc6 : _GEN_1936; // @[control.scala 1315:23 2434:25]
  wire [31:0] _GEN_1946 = 7'h62 == cnt_layer ? 32'h3f521f68 : _GEN_1937; // @[control.scala 1315:23 2435:25]
  wire [7:0] _GEN_1947 = 7'h62 == cnt_layer ? 8'h0 : _GEN_1938; // @[control.scala 1315:23 2436:25]
  wire [31:0] _GEN_1948 = 7'h62 == cnt_layer ? 32'h22b90000 : _GEN_1939; // @[control.scala 1315:23 2437:31]
  wire [31:0] _GEN_1949 = 7'h62 == cnt_layer ? 32'h22d29000 : _GEN_1940; // @[control.scala 1315:23 2438:31]
  wire [15:0] _GEN_1950 = 7'h61 == cnt_layer ? 16'h75fa : _GEN_1941; // @[control.scala 1315:23 2419:25]
  wire [3:0] _GEN_1951 = 7'h61 == cnt_layer ? 4'h8 : _GEN_1942; // @[control.scala 1315:23 2420:25]
  wire [7:0] _GEN_1952 = 7'h61 == cnt_layer ? 8'h4 : _GEN_1943; // @[control.scala 1315:23 2421:25]
  wire [7:0] _GEN_1953 = 7'h61 == cnt_layer ? 8'h4f : _GEN_1944; // @[control.scala 1315:23 2422:25]
  wire [31:0] _GEN_1954 = 7'h61 == cnt_layer ? 32'h3e877e6f : _GEN_1945; // @[control.scala 1315:23 2423:25]
  wire [31:0] _GEN_1955 = 7'h61 == cnt_layer ? 32'h411b4251 : _GEN_1946; // @[control.scala 1315:23 2424:25]
  wire [7:0] _GEN_1956 = 7'h61 == cnt_layer ? 8'h3 : _GEN_1947; // @[control.scala 1315:23 2425:25]
  wire [31:0] _GEN_1957 = 7'h61 == cnt_layer ? 32'h22b48000 : _GEN_1948; // @[control.scala 1315:23 2426:31]
  wire [31:0] _GEN_1958 = 7'h61 == cnt_layer ? 32'h22d28800 : _GEN_1949; // @[control.scala 1315:23 2427:31]
  wire [15:0] _GEN_1959 = 7'h60 == cnt_layer ? 16'h4e42 : _GEN_1950; // @[control.scala 1315:23 2407:25]
  wire [3:0] _GEN_1960 = 7'h60 == cnt_layer ? 4'h7 : _GEN_1951; // @[control.scala 1315:23 2408:25]
  wire [7:0] _GEN_1961 = 7'h60 == cnt_layer ? 8'h0 : _GEN_1952; // @[control.scala 1315:23 2409:25]
  wire [7:0] _GEN_1962 = 7'h60 == cnt_layer ? 8'h74 : _GEN_1953; // @[control.scala 1315:23 2410:25]
  wire [31:0] _GEN_1963 = 7'h60 == cnt_layer ? 32'h3eb2393c : _GEN_1954; // @[control.scala 1315:23 2411:25]
  wire [31:0] _GEN_1964 = 7'h60 == cnt_layer ? 32'h41f78a6d : _GEN_1955; // @[control.scala 1315:23 2412:25]
  wire [7:0] _GEN_1965 = 7'h60 == cnt_layer ? 8'h9 : _GEN_1956; // @[control.scala 1315:23 2413:25]
  wire [31:0] _GEN_1966 = 7'h60 == cnt_layer ? 32'h22b00000 : _GEN_1957; // @[control.scala 1315:23 2414:31]
  wire [31:0] _GEN_1967 = 7'h60 == cnt_layer ? 32'h22d28000 : _GEN_1958; // @[control.scala 1315:23 2415:31]
  wire [15:0] _GEN_1968 = 7'h5f == cnt_layer ? 16'h685b : _GEN_1959; // @[control.scala 1315:23 2396:25]
  wire [3:0] _GEN_1969 = 7'h5f == cnt_layer ? 4'h8 : _GEN_1960; // @[control.scala 1315:23 2397:25]
  wire [7:0] _GEN_1970 = 7'h5f == cnt_layer ? 8'h4 : _GEN_1961; // @[control.scala 1315:23 2398:25]
  wire [7:0] _GEN_1971 = 7'h5f == cnt_layer ? 8'h49 : _GEN_1962; // @[control.scala 1315:23 2399:25]
  wire [31:0] _GEN_1972 = 7'h5f == cnt_layer ? 32'h4003edf4 : _GEN_1963; // @[control.scala 1315:23 2400:25]
  wire [31:0] _GEN_1973 = 7'h5f == cnt_layer ? 32'h3f9063c0 : _GEN_1964; // @[control.scala 1315:23 2401:25]
  wire [7:0] _GEN_1974 = 7'h5f == cnt_layer ? 8'h0 : _GEN_1965; // @[control.scala 1315:23 2402:25]
  wire [31:0] _GEN_1975 = 7'h5f == cnt_layer ? 32'h22a70000 : _GEN_1966; // @[control.scala 1315:23 2403:31]
  wire [31:0] _GEN_1976 = 7'h5f == cnt_layer ? 32'h22d27000 : _GEN_1967; // @[control.scala 1315:23 2404:31]
  wire [15:0] _GEN_1977 = 7'h5e == cnt_layer ? 16'h5539 : _GEN_1968; // @[control.scala 1315:23 2385:25]
  wire [3:0] _GEN_1978 = 7'h5e == cnt_layer ? 4'h8 : _GEN_1969; // @[control.scala 1315:23 2386:25]
  wire [7:0] _GEN_1979 = 7'h5e == cnt_layer ? 8'h4 : _GEN_1970; // @[control.scala 1315:23 2387:25]
  wire [7:0] _GEN_1980 = 7'h5e == cnt_layer ? 8'h50 : _GEN_1971; // @[control.scala 1315:23 2388:25]
  wire [31:0] _GEN_1981 = 7'h5e == cnt_layer ? 32'h3e47b13a : _GEN_1972; // @[control.scala 1315:23 2389:25]
  wire [31:0] _GEN_1982 = 7'h5e == cnt_layer ? 32'h41566442 : _GEN_1973; // @[control.scala 1315:23 2390:25]
  wire [7:0] _GEN_1983 = 7'h5e == cnt_layer ? 8'h4 : _GEN_1974; // @[control.scala 1315:23 2391:25]
  wire [31:0] _GEN_1984 = 7'h5e == cnt_layer ? 32'h22a70000 : _GEN_1975; // @[control.scala 1315:23 2392:31]
  wire [31:0] _GEN_1985 = 7'h5e == cnt_layer ? 32'h22d27000 : _GEN_1976; // @[control.scala 1315:23 2393:31]
  wire [15:0] _GEN_1986 = 7'h5d == cnt_layer ? 16'h6667 : _GEN_1977; // @[control.scala 1315:23 2372:25]
  wire [3:0] _GEN_1987 = 7'h5d == cnt_layer ? 4'h7 : _GEN_1978; // @[control.scala 1315:23 2373:25]
  wire [7:0] _GEN_1988 = 7'h5d == cnt_layer ? 8'h1 : _GEN_1979; // @[control.scala 1315:23 2374:25]
  wire [7:0] _GEN_1989 = 7'h5d == cnt_layer ? 8'h30 : _GEN_1980; // @[control.scala 1315:23 2375:25]
  wire [31:0] _GEN_1990 = 7'h5d == cnt_layer ? 32'h3e3a1e74 : _GEN_1981; // @[control.scala 1315:23 2376:25]
  wire [31:0] _GEN_1991 = 7'h5d == cnt_layer ? 32'h410ad686 : _GEN_1982; // @[control.scala 1315:23 2377:25]
  wire [7:0] _GEN_1992 = 7'h5d == cnt_layer ? 8'h2 : _GEN_1983; // @[control.scala 1315:23 2378:25]
  wire [31:0] _GEN_1993 = 7'h5d == cnt_layer ? 32'h22a28000 : _GEN_1984; // @[control.scala 1315:23 2379:31]
  wire [31:0] _GEN_1994 = 7'h5d == cnt_layer ? 32'h22d26800 : _GEN_1985; // @[control.scala 1315:23 2380:31]
  wire [15:0] _GEN_1995 = 7'h5c == cnt_layer ? 16'h6234 : _GEN_1986; // @[control.scala 1315:23 2361:25]
  wire [3:0] _GEN_1996 = 7'h5c == cnt_layer ? 4'h8 : _GEN_1987; // @[control.scala 1315:23 2362:25]
  wire [7:0] _GEN_1997 = 7'h5c == cnt_layer ? 8'h3 : _GEN_1988; // @[control.scala 1315:23 2363:25]
  wire [7:0] _GEN_1998 = 7'h5c == cnt_layer ? 8'h2d : _GEN_1989; // @[control.scala 1315:23 2364:25]
  wire [31:0] _GEN_1999 = 7'h5c == cnt_layer ? 32'h3f3292ad : _GEN_1990; // @[control.scala 1315:23 2365:25]
  wire [31:0] _GEN_2000 = 7'h5c == cnt_layer ? 32'h400d3592 : _GEN_1991; // @[control.scala 1315:23 2366:25]
  wire [7:0] _GEN_2001 = 7'h5c == cnt_layer ? 8'h1 : _GEN_1992; // @[control.scala 1315:23 2367:25]
  wire [31:0] _GEN_2002 = 7'h5c == cnt_layer ? 32'h229e0000 : _GEN_1993; // @[control.scala 1315:23 2368:31]
  wire [31:0] _GEN_2003 = 7'h5c == cnt_layer ? 32'h22d26000 : _GEN_1994; // @[control.scala 1315:23 2369:31]
  wire [15:0] _GEN_2004 = 7'h5b == cnt_layer ? 16'h643a : _GEN_1995; // @[control.scala 1315:23 2350:25]
  wire [3:0] _GEN_2005 = 7'h5b == cnt_layer ? 4'h8 : _GEN_1996; // @[control.scala 1315:23 2351:25]
  wire [7:0] _GEN_2006 = 7'h5b == cnt_layer ? 8'h3 : _GEN_1997; // @[control.scala 1315:23 2352:25]
  wire [7:0] _GEN_2007 = 7'h5b == cnt_layer ? 8'h4e : _GEN_1998; // @[control.scala 1315:23 2353:25]
  wire [31:0] _GEN_2008 = 7'h5b == cnt_layer ? 32'h3e90adec : _GEN_1999; // @[control.scala 1315:23 2354:25]
  wire [31:0] _GEN_2009 = 7'h5b == cnt_layer ? 32'h41103fe0 : _GEN_2000; // @[control.scala 1315:23 2355:25]
  wire [7:0] _GEN_2010 = 7'h5b == cnt_layer ? 8'h3 : _GEN_2001; // @[control.scala 1315:23 2356:25]
  wire [31:0] _GEN_2011 = 7'h5b == cnt_layer ? 32'h22998000 : _GEN_2002; // @[control.scala 1315:23 2357:31]
  wire [31:0] _GEN_2012 = 7'h5b == cnt_layer ? 32'h22d25800 : _GEN_2003; // @[control.scala 1315:23 2358:31]
  wire [15:0] _GEN_2013 = 7'h5a == cnt_layer ? 16'h56ee : _GEN_2004; // @[control.scala 1315:23 2338:25]
  wire [3:0] _GEN_2014 = 7'h5a == cnt_layer ? 4'h7 : _GEN_2005; // @[control.scala 1315:23 2339:25]
  wire [7:0] _GEN_2015 = 7'h5a == cnt_layer ? 8'h1 : _GEN_2006; // @[control.scala 1315:23 2340:25]
  wire [7:0] _GEN_2016 = 7'h5a == cnt_layer ? 8'h32 : _GEN_2007; // @[control.scala 1315:23 2341:25]
  wire [31:0] _GEN_2017 = 7'h5a == cnt_layer ? 32'h3e69ed97 : _GEN_2008; // @[control.scala 1315:23 2342:25]
  wire [31:0] _GEN_2018 = 7'h5a == cnt_layer ? 32'h40e4d2b1 : _GEN_2009; // @[control.scala 1315:23 2343:25]
  wire [7:0] _GEN_2019 = 7'h5a == cnt_layer ? 8'h2 : _GEN_2010; // @[control.scala 1315:23 2344:25]
  wire [31:0] _GEN_2020 = 7'h5a == cnt_layer ? 32'h22950000 : _GEN_2011; // @[control.scala 1315:23 2345:31]
  wire [31:0] _GEN_2021 = 7'h5a == cnt_layer ? 32'h22d25000 : _GEN_2012; // @[control.scala 1315:23 2346:31]
  wire [15:0] _GEN_2022 = 7'h59 == cnt_layer ? 16'h516d : _GEN_2013; // @[control.scala 1315:23 2327:25]
  wire [3:0] _GEN_2023 = 7'h59 == cnt_layer ? 4'h7 : _GEN_2014; // @[control.scala 1315:23 2328:25]
  wire [7:0] _GEN_2024 = 7'h59 == cnt_layer ? 8'h2 : _GEN_2015; // @[control.scala 1315:23 2329:25]
  wire [7:0] _GEN_2025 = 7'h59 == cnt_layer ? 8'h31 : _GEN_2016; // @[control.scala 1315:23 2330:25]
  wire [31:0] _GEN_2026 = 7'h59 == cnt_layer ? 32'h3f403ce5 : _GEN_2017; // @[control.scala 1315:23 2331:25]
  wire [31:0] _GEN_2027 = 7'h59 == cnt_layer ? 32'h400a35e8 : _GEN_2018; // @[control.scala 1315:23 2332:25]
  wire [7:0] _GEN_2028 = 7'h59 == cnt_layer ? 8'h1 : _GEN_2019; // @[control.scala 1315:23 2333:25]
  wire [31:0] _GEN_2029 = 7'h59 == cnt_layer ? 32'h22908000 : _GEN_2020; // @[control.scala 1315:23 2334:31]
  wire [31:0] _GEN_2030 = 7'h59 == cnt_layer ? 32'h22d24800 : _GEN_2021; // @[control.scala 1315:23 2335:31]
  wire [15:0] _GEN_2031 = 7'h58 == cnt_layer ? 16'h6968 : _GEN_2022; // @[control.scala 1315:23 2316:25]
  wire [3:0] _GEN_2032 = 7'h58 == cnt_layer ? 4'h8 : _GEN_2023; // @[control.scala 1315:23 2317:25]
  wire [7:0] _GEN_2033 = 7'h58 == cnt_layer ? 8'h4 : _GEN_2024; // @[control.scala 1315:23 2318:25]
  wire [7:0] _GEN_2034 = 7'h58 == cnt_layer ? 8'h4c : _GEN_2025; // @[control.scala 1315:23 2319:25]
  wire [31:0] _GEN_2035 = 7'h58 == cnt_layer ? 32'h3e9f26a6 : _GEN_2026; // @[control.scala 1315:23 2320:25]
  wire [31:0] _GEN_2036 = 7'h58 == cnt_layer ? 32'h40fa153b : _GEN_2027; // @[control.scala 1315:23 2321:25]
  wire [7:0] _GEN_2037 = 7'h58 == cnt_layer ? 8'h2 : _GEN_2028; // @[control.scala 1315:23 2322:25]
  wire [31:0] _GEN_2038 = 7'h58 == cnt_layer ? 32'h228c0000 : _GEN_2029; // @[control.scala 1315:23 2323:31]
  wire [31:0] _GEN_2039 = 7'h58 == cnt_layer ? 32'h22d24000 : _GEN_2030; // @[control.scala 1315:23 2324:31]
  wire [15:0] _GEN_2040 = 7'h57 == cnt_layer ? 16'h6bb4 : _GEN_2031; // @[control.scala 1315:23 2304:25]
  wire [3:0] _GEN_2041 = 7'h57 == cnt_layer ? 4'h8 : _GEN_2032; // @[control.scala 1315:23 2305:25]
  wire [7:0] _GEN_2042 = 7'h57 == cnt_layer ? 8'h1 : _GEN_2033; // @[control.scala 1315:23 2306:25]
  wire [7:0] _GEN_2043 = 7'h57 == cnt_layer ? 8'h20 : _GEN_2034; // @[control.scala 1315:23 2307:25]
  wire [31:0] _GEN_2044 = 7'h57 == cnt_layer ? 32'h3e9d496f : _GEN_2035; // @[control.scala 1315:23 2308:25]
  wire [31:0] _GEN_2045 = 7'h57 == cnt_layer ? 32'h408a58c4 : _GEN_2036; // @[control.scala 1315:23 2309:25]
  wire [7:0] _GEN_2046 = 7'h57 == cnt_layer ? 8'h1 : _GEN_2037; // @[control.scala 1315:23 2310:25]
  wire [31:0] _GEN_2047 = 7'h57 == cnt_layer ? 32'h22878000 : _GEN_2038; // @[control.scala 1315:23 2311:31]
  wire [31:0] _GEN_2048 = 7'h57 == cnt_layer ? 32'h22d23800 : _GEN_2039; // @[control.scala 1315:23 2312:31]
  wire [15:0] _GEN_2049 = 7'h56 == cnt_layer ? 16'h4f34 : _GEN_2040; // @[control.scala 1315:23 2293:25]
  wire [3:0] _GEN_2050 = 7'h56 == cnt_layer ? 4'h7 : _GEN_2041; // @[control.scala 1315:23 2294:25]
  wire [7:0] _GEN_2051 = 7'h56 == cnt_layer ? 8'h4 : _GEN_2042; // @[control.scala 1315:23 2295:25]
  wire [7:0] _GEN_2052 = 7'h56 == cnt_layer ? 8'h35 : _GEN_2043; // @[control.scala 1315:23 2296:25]
  wire [31:0] _GEN_2053 = 7'h56 == cnt_layer ? 32'h3f367e4b : _GEN_2044; // @[control.scala 1315:23 2297:25]
  wire [31:0] _GEN_2054 = 7'h56 == cnt_layer ? 32'h401987b7 : _GEN_2045; // @[control.scala 1315:23 2298:25]
  wire [7:0] _GEN_2055 = 7'h56 == cnt_layer ? 8'h1 : _GEN_2046; // @[control.scala 1315:23 2299:25]
  wire [31:0] _GEN_2056 = 7'h56 == cnt_layer ? 32'h22830000 : _GEN_2047; // @[control.scala 1315:23 2300:31]
  wire [31:0] _GEN_2057 = 7'h56 == cnt_layer ? 32'h22d23000 : _GEN_2048; // @[control.scala 1315:23 2301:31]
  wire [15:0] _GEN_2058 = 7'h55 == cnt_layer ? 16'h565d : _GEN_2049; // @[control.scala 1315:23 2282:25]
  wire [3:0] _GEN_2059 = 7'h55 == cnt_layer ? 4'h8 : _GEN_2050; // @[control.scala 1315:23 2283:25]
  wire [7:0] _GEN_2060 = 7'h55 == cnt_layer ? 8'h4 : _GEN_2051; // @[control.scala 1315:23 2284:25]
  wire [7:0] _GEN_2061 = 7'h55 == cnt_layer ? 8'h55 : _GEN_2052; // @[control.scala 1315:23 2285:25]
  wire [31:0] _GEN_2062 = 7'h55 == cnt_layer ? 32'h3e6dc373 : _GEN_2053; // @[control.scala 1315:23 2286:25]
  wire [31:0] _GEN_2063 = 7'h55 == cnt_layer ? 32'h414b81af : _GEN_2054; // @[control.scala 1315:23 2287:25]
  wire [7:0] _GEN_2064 = 7'h55 == cnt_layer ? 8'h4 : _GEN_2055; // @[control.scala 1315:23 2288:25]
  wire [31:0] _GEN_2065 = 7'h55 == cnt_layer ? 32'h227e8000 : _GEN_2056; // @[control.scala 1315:23 2289:31]
  wire [31:0] _GEN_2066 = 7'h55 == cnt_layer ? 32'h22d22800 : _GEN_2057; // @[control.scala 1315:23 2290:31]
  wire [15:0] _GEN_2067 = 7'h54 == cnt_layer ? 16'h67a3 : _GEN_2058; // @[control.scala 1315:23 2269:25]
  wire [3:0] _GEN_2068 = 7'h54 == cnt_layer ? 4'h7 : _GEN_2059; // @[control.scala 1315:23 2270:25]
  wire [7:0] _GEN_2069 = 7'h54 == cnt_layer ? 8'h2 : _GEN_2060; // @[control.scala 1315:23 2271:25]
  wire [7:0] _GEN_2070 = 7'h54 == cnt_layer ? 8'h5b : _GEN_2061; // @[control.scala 1315:23 2272:25]
  wire [31:0] _GEN_2071 = 7'h54 == cnt_layer ? 32'h3eb5a49f : _GEN_2062; // @[control.scala 1315:23 2273:25]
  wire [31:0] _GEN_2072 = 7'h54 == cnt_layer ? 32'h411dc0a1 : _GEN_2063; // @[control.scala 1315:23 2274:25]
  wire [7:0] _GEN_2073 = 7'h54 == cnt_layer ? 8'h3 : _GEN_2064; // @[control.scala 1315:23 2275:25]
  wire [31:0] _GEN_2074 = 7'h54 == cnt_layer ? 32'h227a0000 : _GEN_2065; // @[control.scala 1315:23 2276:31]
  wire [31:0] _GEN_2075 = 7'h54 == cnt_layer ? 32'h22d22000 : _GEN_2066; // @[control.scala 1315:23 2277:31]
  wire [15:0] _GEN_2076 = 7'h53 == cnt_layer ? 16'h1 : _GEN_2067; // @[control.scala 1315:23 2258:25]
  wire [3:0] _GEN_2077 = 7'h53 == cnt_layer ? 4'h0 : _GEN_2068; // @[control.scala 1315:23 2259:25]
  wire [7:0] _GEN_2078 = 7'h53 == cnt_layer ? 8'h0 : _GEN_2069; // @[control.scala 1315:23 2260:25]
  wire [7:0] _GEN_2079 = 7'h53 == cnt_layer ? 8'h0 : _GEN_2070; // @[control.scala 1315:23 2261:25]
  wire [31:0] _GEN_2080 = 7'h53 == cnt_layer ? 32'h3f800000 : _GEN_2071; // @[control.scala 1315:23 2262:25]
  wire [31:0] _GEN_2081 = 7'h53 == cnt_layer ? 32'h3f800000 : _GEN_2072; // @[control.scala 1315:23 2263:25]
  wire [7:0] _GEN_2082 = 7'h53 == cnt_layer ? 8'h0 : _GEN_2073; // @[control.scala 1315:23 2264:25]
  wire [31:0] _GEN_2083 = 7'h53 == cnt_layer ? 32'h22758000 : _GEN_2074; // @[control.scala 1315:23 2265:31]
  wire [31:0] _GEN_2084 = 7'h53 == cnt_layer ? 32'h22d21800 : _GEN_2075; // @[control.scala 1315:23 2266:31]
  wire [15:0] _GEN_2085 = 7'h52 == cnt_layer ? 16'h1 : _GEN_2076; // @[control.scala 1315:23 2247:25]
  wire [3:0] _GEN_2086 = 7'h52 == cnt_layer ? 4'h0 : _GEN_2077; // @[control.scala 1315:23 2248:25]
  wire [7:0] _GEN_2087 = 7'h52 == cnt_layer ? 8'h0 : _GEN_2078; // @[control.scala 1315:23 2249:25]
  wire [7:0] _GEN_2088 = 7'h52 == cnt_layer ? 8'h0 : _GEN_2079; // @[control.scala 1315:23 2250:25]
  wire [31:0] _GEN_2089 = 7'h52 == cnt_layer ? 32'h3f800000 : _GEN_2080; // @[control.scala 1315:23 2251:25]
  wire [31:0] _GEN_2090 = 7'h52 == cnt_layer ? 32'h3f800000 : _GEN_2081; // @[control.scala 1315:23 2252:25]
  wire [7:0] _GEN_2091 = 7'h52 == cnt_layer ? 8'h0 : _GEN_2082; // @[control.scala 1315:23 2253:25]
  wire [31:0] _GEN_2092 = 7'h52 == cnt_layer ? 32'h22710000 : _GEN_2083; // @[control.scala 1315:23 2254:31]
  wire [31:0] _GEN_2093 = 7'h52 == cnt_layer ? 32'h22d21000 : _GEN_2084; // @[control.scala 1315:23 2255:31]
  wire [15:0] _GEN_2094 = 7'h51 == cnt_layer ? 16'h1 : _GEN_2085; // @[control.scala 1315:23 2236:25]
  wire [3:0] _GEN_2095 = 7'h51 == cnt_layer ? 4'h0 : _GEN_2086; // @[control.scala 1315:23 2237:25]
  wire [7:0] _GEN_2096 = 7'h51 == cnt_layer ? 8'h0 : _GEN_2087; // @[control.scala 1315:23 2238:25]
  wire [7:0] _GEN_2097 = 7'h51 == cnt_layer ? 8'h0 : _GEN_2088; // @[control.scala 1315:23 2239:25]
  wire [31:0] _GEN_2098 = 7'h51 == cnt_layer ? 32'h3f800000 : _GEN_2089; // @[control.scala 1315:23 2240:25]
  wire [31:0] _GEN_2099 = 7'h51 == cnt_layer ? 32'h3f800000 : _GEN_2090; // @[control.scala 1315:23 2241:25]
  wire [7:0] _GEN_2100 = 7'h51 == cnt_layer ? 8'h0 : _GEN_2091; // @[control.scala 1315:23 2242:25]
  wire [31:0] _GEN_2101 = 7'h51 == cnt_layer ? 32'h226c8000 : _GEN_2092; // @[control.scala 1315:23 2243:31]
  wire [31:0] _GEN_2102 = 7'h51 == cnt_layer ? 32'h22d20800 : _GEN_2093; // @[control.scala 1315:23 2244:31]
  wire [15:0] _GEN_2103 = 7'h50 == cnt_layer ? 16'h1 : _GEN_2094; // @[control.scala 1315:23 2225:25]
  wire [3:0] _GEN_2104 = 7'h50 == cnt_layer ? 4'h0 : _GEN_2095; // @[control.scala 1315:23 2226:25]
  wire [7:0] _GEN_2105 = 7'h50 == cnt_layer ? 8'h0 : _GEN_2096; // @[control.scala 1315:23 2227:25]
  wire [7:0] _GEN_2106 = 7'h50 == cnt_layer ? 8'h0 : _GEN_2097; // @[control.scala 1315:23 2228:25]
  wire [31:0] _GEN_2107 = 7'h50 == cnt_layer ? 32'h3f800000 : _GEN_2098; // @[control.scala 1315:23 2229:25]
  wire [31:0] _GEN_2108 = 7'h50 == cnt_layer ? 32'h3f800000 : _GEN_2099; // @[control.scala 1315:23 2230:25]
  wire [7:0] _GEN_2109 = 7'h50 == cnt_layer ? 8'h0 : _GEN_2100; // @[control.scala 1315:23 2231:25]
  wire [31:0] _GEN_2110 = 7'h50 == cnt_layer ? 32'h22680000 : _GEN_2101; // @[control.scala 1315:23 2232:31]
  wire [31:0] _GEN_2111 = 7'h50 == cnt_layer ? 32'h22d20000 : _GEN_2102; // @[control.scala 1315:23 2233:31]
  wire [15:0] _GEN_2112 = 7'h4f == cnt_layer ? 16'h45f1 : _GEN_2103; // @[control.scala 1315:23 2214:25]
  wire [3:0] _GEN_2113 = 7'h4f == cnt_layer ? 4'h7 : _GEN_2104; // @[control.scala 1315:23 2215:25]
  wire [7:0] _GEN_2114 = 7'h4f == cnt_layer ? 8'h4 : _GEN_2105; // @[control.scala 1315:23 2216:25]
  wire [7:0] _GEN_2115 = 7'h4f == cnt_layer ? 8'h3e : _GEN_2106; // @[control.scala 1315:23 2217:25]
  wire [31:0] _GEN_2116 = 7'h4f == cnt_layer ? 32'h3e730a55 : _GEN_2107; // @[control.scala 1315:23 2218:25]
  wire [31:0] _GEN_2117 = 7'h4f == cnt_layer ? 32'h41018c19 : _GEN_2108; // @[control.scala 1315:23 2219:25]
  wire [7:0] _GEN_2118 = 7'h4f == cnt_layer ? 8'h2 : _GEN_2109; // @[control.scala 1315:23 2220:25]
  wire [31:0] _GEN_2119 = 7'h4f == cnt_layer ? 32'h22638000 : _GEN_2110; // @[control.scala 1315:23 2221:31]
  wire [31:0] _GEN_2120 = 7'h4f == cnt_layer ? 32'h22d1f800 : _GEN_2111; // @[control.scala 1315:23 2222:31]
  wire [15:0] _GEN_2121 = 7'h4e == cnt_layer ? 16'h426e : _GEN_2112; // @[control.scala 1315:23 2203:25]
  wire [3:0] _GEN_2122 = 7'h4e == cnt_layer ? 4'h7 : _GEN_2113; // @[control.scala 1315:23 2204:25]
  wire [7:0] _GEN_2123 = 7'h4e == cnt_layer ? 8'h3 : _GEN_2114; // @[control.scala 1315:23 2205:25]
  wire [7:0] _GEN_2124 = 7'h4e == cnt_layer ? 8'h49 : _GEN_2115; // @[control.scala 1315:23 2206:25]
  wire [31:0] _GEN_2125 = 7'h4e == cnt_layer ? 32'h3e2afdfc : _GEN_2116; // @[control.scala 1315:23 2207:25]
  wire [31:0] _GEN_2126 = 7'h4e == cnt_layer ? 32'h4158ffd1 : _GEN_2117; // @[control.scala 1315:23 2208:25]
  wire [7:0] _GEN_2127 = 7'h4e == cnt_layer ? 8'h4 : _GEN_2118; // @[control.scala 1315:23 2209:25]
  wire [31:0] _GEN_2128 = 7'h4e == cnt_layer ? 32'h225f0000 : _GEN_2119; // @[control.scala 1315:23 2210:31]
  wire [31:0] _GEN_2129 = 7'h4e == cnt_layer ? 32'h22d1f000 : _GEN_2120; // @[control.scala 1315:23 2211:31]
  wire [15:0] _GEN_2130 = 7'h4d == cnt_layer ? 16'h5edf : _GEN_2121; // @[control.scala 1315:23 2192:25]
  wire [3:0] _GEN_2131 = 7'h4d == cnt_layer ? 4'h7 : _GEN_2122; // @[control.scala 1315:23 2193:25]
  wire [7:0] _GEN_2132 = 7'h4d == cnt_layer ? 8'h3 : _GEN_2123; // @[control.scala 1315:23 2194:25]
  wire [7:0] _GEN_2133 = 7'h4d == cnt_layer ? 8'h45 : _GEN_2124; // @[control.scala 1315:23 2195:25]
  wire [31:0] _GEN_2134 = 7'h4d == cnt_layer ? 32'h3e618f3a : _GEN_2125; // @[control.scala 1315:23 2196:25]
  wire [31:0] _GEN_2135 = 7'h4d == cnt_layer ? 32'h411bc576 : _GEN_2126; // @[control.scala 1315:23 2197:25]
  wire [7:0] _GEN_2136 = 7'h4d == cnt_layer ? 8'h3 : _GEN_2127; // @[control.scala 1315:23 2198:25]
  wire [31:0] _GEN_2137 = 7'h4d == cnt_layer ? 32'h225a8000 : _GEN_2128; // @[control.scala 1315:23 2199:31]
  wire [31:0] _GEN_2138 = 7'h4d == cnt_layer ? 32'h22d1e800 : _GEN_2129; // @[control.scala 1315:23 2200:31]
  wire [15:0] _GEN_2139 = 7'h4c == cnt_layer ? 16'h48b2 : _GEN_2130; // @[control.scala 1315:23 2179:25]
  wire [3:0] _GEN_2140 = 7'h4c == cnt_layer ? 4'h9 : _GEN_2131; // @[control.scala 1315:23 2180:25]
  wire [7:0] _GEN_2141 = 7'h4c == cnt_layer ? 8'h4 : _GEN_2132; // @[control.scala 1315:23 2181:25]
  wire [7:0] _GEN_2142 = 7'h4c == cnt_layer ? 8'h41 : _GEN_2133; // @[control.scala 1315:23 2182:25]
  wire [31:0] _GEN_2143 = 7'h4c == cnt_layer ? 32'h3e59a081 : _GEN_2134; // @[control.scala 1315:23 2183:25]
  wire [31:0] _GEN_2144 = 7'h4c == cnt_layer ? 32'h4116289a : _GEN_2135; // @[control.scala 1315:23 2184:25]
  wire [7:0] _GEN_2145 = 7'h4c == cnt_layer ? 8'h3 : _GEN_2136; // @[control.scala 1315:23 2185:25]
  wire [31:0] _GEN_2146 = 7'h4c == cnt_layer ? 32'h22560000 : _GEN_2137; // @[control.scala 1315:23 2186:31]
  wire [31:0] _GEN_2147 = 7'h4c == cnt_layer ? 32'h22d1e000 : _GEN_2138; // @[control.scala 1315:23 2187:31]
  wire [15:0] _GEN_2148 = 7'h4b == cnt_layer ? 16'h6fe9 : _GEN_2139; // @[control.scala 1315:23 2167:25]
  wire [3:0] _GEN_2149 = 7'h4b == cnt_layer ? 4'h7 : _GEN_2140; // @[control.scala 1315:23 2168:25]
  wire [7:0] _GEN_2150 = 7'h4b == cnt_layer ? 8'h3 : _GEN_2141; // @[control.scala 1315:23 2169:25]
  wire [7:0] _GEN_2151 = 7'h4b == cnt_layer ? 8'h58 : _GEN_2142; // @[control.scala 1315:23 2170:25]
  wire [31:0] _GEN_2152 = 7'h4b == cnt_layer ? 32'h3e4d4e93 : _GEN_2143; // @[control.scala 1315:23 2171:25]
  wire [31:0] _GEN_2153 = 7'h4b == cnt_layer ? 32'h417a3158 : _GEN_2144; // @[control.scala 1315:23 2172:25]
  wire [7:0] _GEN_2154 = 7'h4b == cnt_layer ? 8'h4 : _GEN_2145; // @[control.scala 1315:23 2173:25]
  wire [31:0] _GEN_2155 = 7'h4b == cnt_layer ? 32'h22518000 : _GEN_2146; // @[control.scala 1315:23 2174:31]
  wire [31:0] _GEN_2156 = 7'h4b == cnt_layer ? 32'h22d1d800 : _GEN_2147; // @[control.scala 1315:23 2175:31]
  wire [15:0] _GEN_2157 = 7'h4a == cnt_layer ? 16'h1 : _GEN_2148; // @[control.scala 1315:23 2156:25]
  wire [3:0] _GEN_2158 = 7'h4a == cnt_layer ? 4'h0 : _GEN_2149; // @[control.scala 1315:23 2157:25]
  wire [7:0] _GEN_2159 = 7'h4a == cnt_layer ? 8'h0 : _GEN_2150; // @[control.scala 1315:23 2158:25]
  wire [7:0] _GEN_2160 = 7'h4a == cnt_layer ? 8'h0 : _GEN_2151; // @[control.scala 1315:23 2159:25]
  wire [31:0] _GEN_2161 = 7'h4a == cnt_layer ? 32'h3f800000 : _GEN_2152; // @[control.scala 1315:23 2160:25]
  wire [31:0] _GEN_2162 = 7'h4a == cnt_layer ? 32'h3f800000 : _GEN_2153; // @[control.scala 1315:23 2161:25]
  wire [7:0] _GEN_2163 = 7'h4a == cnt_layer ? 8'h0 : _GEN_2154; // @[control.scala 1315:23 2162:25]
  wire [31:0] _GEN_2164 = 7'h4a == cnt_layer ? 32'h224d0000 : _GEN_2155; // @[control.scala 1315:23 2163:31]
  wire [31:0] _GEN_2165 = 7'h4a == cnt_layer ? 32'h22d1d000 : _GEN_2156; // @[control.scala 1315:23 2164:31]
  wire [15:0] _GEN_2166 = 7'h49 == cnt_layer ? 16'h1 : _GEN_2157; // @[control.scala 1315:23 2145:25]
  wire [3:0] _GEN_2167 = 7'h49 == cnt_layer ? 4'h0 : _GEN_2158; // @[control.scala 1315:23 2146:25]
  wire [7:0] _GEN_2168 = 7'h49 == cnt_layer ? 8'h0 : _GEN_2159; // @[control.scala 1315:23 2147:25]
  wire [7:0] _GEN_2169 = 7'h49 == cnt_layer ? 8'h0 : _GEN_2160; // @[control.scala 1315:23 2148:25]
  wire [31:0] _GEN_2170 = 7'h49 == cnt_layer ? 32'h3f800000 : _GEN_2161; // @[control.scala 1315:23 2149:25]
  wire [31:0] _GEN_2171 = 7'h49 == cnt_layer ? 32'h3f800000 : _GEN_2162; // @[control.scala 1315:23 2150:25]
  wire [7:0] _GEN_2172 = 7'h49 == cnt_layer ? 8'h0 : _GEN_2163; // @[control.scala 1315:23 2151:25]
  wire [31:0] _GEN_2173 = 7'h49 == cnt_layer ? 32'h22488000 : _GEN_2164; // @[control.scala 1315:23 2152:31]
  wire [31:0] _GEN_2174 = 7'h49 == cnt_layer ? 32'h22d1c800 : _GEN_2165; // @[control.scala 1315:23 2153:31]
  wire [15:0] _GEN_2175 = 7'h48 == cnt_layer ? 16'h1 : _GEN_2166; // @[control.scala 1315:23 2134:25]
  wire [3:0] _GEN_2176 = 7'h48 == cnt_layer ? 4'h0 : _GEN_2167; // @[control.scala 1315:23 2135:25]
  wire [7:0] _GEN_2177 = 7'h48 == cnt_layer ? 8'h0 : _GEN_2168; // @[control.scala 1315:23 2136:25]
  wire [7:0] _GEN_2178 = 7'h48 == cnt_layer ? 8'h0 : _GEN_2169; // @[control.scala 1315:23 2137:25]
  wire [31:0] _GEN_2179 = 7'h48 == cnt_layer ? 32'h3f800000 : _GEN_2170; // @[control.scala 1315:23 2138:25]
  wire [31:0] _GEN_2180 = 7'h48 == cnt_layer ? 32'h3f800000 : _GEN_2171; // @[control.scala 1315:23 2139:25]
  wire [7:0] _GEN_2181 = 7'h48 == cnt_layer ? 8'h0 : _GEN_2172; // @[control.scala 1315:23 2140:25]
  wire [31:0] _GEN_2182 = 7'h48 == cnt_layer ? 32'h22440000 : _GEN_2173; // @[control.scala 1315:23 2141:31]
  wire [31:0] _GEN_2183 = 7'h48 == cnt_layer ? 32'h22d1c000 : _GEN_2174; // @[control.scala 1315:23 2142:31]
  wire [15:0] _GEN_2184 = 7'h47 == cnt_layer ? 16'h1 : _GEN_2175; // @[control.scala 1315:23 2123:25]
  wire [3:0] _GEN_2185 = 7'h47 == cnt_layer ? 4'h0 : _GEN_2176; // @[control.scala 1315:23 2124:25]
  wire [7:0] _GEN_2186 = 7'h47 == cnt_layer ? 8'h0 : _GEN_2177; // @[control.scala 1315:23 2125:25]
  wire [7:0] _GEN_2187 = 7'h47 == cnt_layer ? 8'h0 : _GEN_2178; // @[control.scala 1315:23 2126:25]
  wire [31:0] _GEN_2188 = 7'h47 == cnt_layer ? 32'h3f800000 : _GEN_2179; // @[control.scala 1315:23 2127:25]
  wire [31:0] _GEN_2189 = 7'h47 == cnt_layer ? 32'h3f800000 : _GEN_2180; // @[control.scala 1315:23 2128:25]
  wire [7:0] _GEN_2190 = 7'h47 == cnt_layer ? 8'h0 : _GEN_2181; // @[control.scala 1315:23 2129:25]
  wire [31:0] _GEN_2191 = 7'h47 == cnt_layer ? 32'h223f8000 : _GEN_2182; // @[control.scala 1315:23 2130:31]
  wire [31:0] _GEN_2192 = 7'h47 == cnt_layer ? 32'h22d1b800 : _GEN_2183; // @[control.scala 1315:23 2131:31]
  wire [15:0] _GEN_2193 = 7'h46 == cnt_layer ? 16'h755c : _GEN_2184; // @[control.scala 1315:23 2112:25]
  wire [3:0] _GEN_2194 = 7'h46 == cnt_layer ? 4'h8 : _GEN_2185; // @[control.scala 1315:23 2113:25]
  wire [7:0] _GEN_2195 = 7'h46 == cnt_layer ? 8'h6 : _GEN_2186; // @[control.scala 1315:23 2114:25]
  wire [7:0] _GEN_2196 = 7'h46 == cnt_layer ? 8'h47 : _GEN_2187; // @[control.scala 1315:23 2115:25]
  wire [31:0] _GEN_2197 = 7'h46 == cnt_layer ? 32'h3e6c4438 : _GEN_2188; // @[control.scala 1315:23 2116:25]
  wire [31:0] _GEN_2198 = 7'h46 == cnt_layer ? 32'h41192dca : _GEN_2189; // @[control.scala 1315:23 2117:25]
  wire [7:0] _GEN_2199 = 7'h46 == cnt_layer ? 8'h3 : _GEN_2190; // @[control.scala 1315:23 2118:25]
  wire [31:0] _GEN_2200 = 7'h46 == cnt_layer ? 32'h223b0000 : _GEN_2191; // @[control.scala 1315:23 2119:31]
  wire [31:0] _GEN_2201 = 7'h46 == cnt_layer ? 32'h22d1b000 : _GEN_2192; // @[control.scala 1315:23 2120:31]
  wire [15:0] _GEN_2202 = 7'h45 == cnt_layer ? 16'h450e : _GEN_2193; // @[control.scala 1315:23 2101:25]
  wire [3:0] _GEN_2203 = 7'h45 == cnt_layer ? 4'h7 : _GEN_2194; // @[control.scala 1315:23 2102:25]
  wire [7:0] _GEN_2204 = 7'h45 == cnt_layer ? 8'h3 : _GEN_2195; // @[control.scala 1315:23 2103:25]
  wire [7:0] _GEN_2205 = 7'h45 == cnt_layer ? 8'h50 : _GEN_2196; // @[control.scala 1315:23 2104:25]
  wire [31:0] _GEN_2206 = 7'h45 == cnt_layer ? 32'h3df96b8d : _GEN_2197; // @[control.scala 1315:23 2105:25]
  wire [31:0] _GEN_2207 = 7'h45 == cnt_layer ? 32'h41a8a6f9 : _GEN_2198; // @[control.scala 1315:23 2106:25]
  wire [7:0] _GEN_2208 = 7'h45 == cnt_layer ? 8'h6 : _GEN_2199; // @[control.scala 1315:23 2107:25]
  wire [31:0] _GEN_2209 = 7'h45 == cnt_layer ? 32'h22368000 : _GEN_2200; // @[control.scala 1315:23 2108:31]
  wire [31:0] _GEN_2210 = 7'h45 == cnt_layer ? 32'h22d1a800 : _GEN_2201; // @[control.scala 1315:23 2109:31]
  wire [15:0] _GEN_2211 = 7'h44 == cnt_layer ? 16'h697d : _GEN_2202; // @[control.scala 1315:23 2090:25]
  wire [3:0] _GEN_2212 = 7'h44 == cnt_layer ? 4'h8 : _GEN_2203; // @[control.scala 1315:23 2091:25]
  wire [7:0] _GEN_2213 = 7'h44 == cnt_layer ? 8'h4 : _GEN_2204; // @[control.scala 1315:23 2092:25]
  wire [7:0] _GEN_2214 = 7'h44 == cnt_layer ? 8'h44 : _GEN_2205; // @[control.scala 1315:23 2093:25]
  wire [31:0] _GEN_2215 = 7'h44 == cnt_layer ? 32'h3e418575 : _GEN_2206; // @[control.scala 1315:23 2094:25]
  wire [31:0] _GEN_2216 = 7'h44 == cnt_layer ? 32'h41325df1 : _GEN_2207; // @[control.scala 1315:23 2095:25]
  wire [7:0] _GEN_2217 = 7'h44 == cnt_layer ? 8'h3 : _GEN_2208; // @[control.scala 1315:23 2096:25]
  wire [31:0] _GEN_2218 = 7'h44 == cnt_layer ? 32'h22320000 : _GEN_2209; // @[control.scala 1315:23 2097:31]
  wire [31:0] _GEN_2219 = 7'h44 == cnt_layer ? 32'h22d1a000 : _GEN_2210; // @[control.scala 1315:23 2098:31]
  wire [15:0] _GEN_2220 = 7'h43 == cnt_layer ? 16'h5517 : _GEN_2211; // @[control.scala 1315:23 2077:25]
  wire [3:0] _GEN_2221 = 7'h43 == cnt_layer ? 4'h8 : _GEN_2212; // @[control.scala 1315:23 2078:25]
  wire [7:0] _GEN_2222 = 7'h43 == cnt_layer ? 8'h4 : _GEN_2213; // @[control.scala 1315:23 2079:25]
  wire [7:0] _GEN_2223 = 7'h43 == cnt_layer ? 8'h46 : _GEN_2214; // @[control.scala 1315:23 2080:25]
  wire [31:0] _GEN_2224 = 7'h43 == cnt_layer ? 32'h3e19caee : _GEN_2215; // @[control.scala 1315:23 2081:25]
  wire [31:0] _GEN_2225 = 7'h43 == cnt_layer ? 32'h41678464 : _GEN_2216; // @[control.scala 1315:23 2082:25]
  wire [7:0] _GEN_2226 = 7'h43 == cnt_layer ? 8'h4 : _GEN_2217; // @[control.scala 1315:23 2083:25]
  wire [31:0] _GEN_2227 = 7'h43 == cnt_layer ? 32'h222d8000 : _GEN_2218; // @[control.scala 1315:23 2084:31]
  wire [31:0] _GEN_2228 = 7'h43 == cnt_layer ? 32'h22d19800 : _GEN_2219; // @[control.scala 1315:23 2085:31]
  wire [15:0] _GEN_2229 = 7'h42 == cnt_layer ? 16'h4745 : _GEN_2220; // @[control.scala 1315:23 2065:25]
  wire [3:0] _GEN_2230 = 7'h42 == cnt_layer ? 4'h7 : _GEN_2221; // @[control.scala 1315:23 2066:25]
  wire [7:0] _GEN_2231 = 7'h42 == cnt_layer ? 8'h4 : _GEN_2222; // @[control.scala 1315:23 2067:25]
  wire [7:0] _GEN_2232 = 7'h42 == cnt_layer ? 8'h4b : _GEN_2223; // @[control.scala 1315:23 2068:25]
  wire [31:0] _GEN_2233 = 7'h42 == cnt_layer ? 32'h3e1e8114 : _GEN_2224; // @[control.scala 1315:23 2069:25]
  wire [31:0] _GEN_2234 = 7'h42 == cnt_layer ? 32'h4173e8bc : _GEN_2225; // @[control.scala 1315:23 2070:25]
  wire [7:0] _GEN_2235 = 7'h42 == cnt_layer ? 8'h4 : _GEN_2226; // @[control.scala 1315:23 2071:25]
  wire [31:0] _GEN_2236 = 7'h42 == cnt_layer ? 32'h22290000 : _GEN_2227; // @[control.scala 1315:23 2072:31]
  wire [31:0] _GEN_2237 = 7'h42 == cnt_layer ? 32'h22d19000 : _GEN_2228; // @[control.scala 1315:23 2073:31]
  wire [15:0] _GEN_2238 = 7'h41 == cnt_layer ? 16'h1 : _GEN_2229; // @[control.scala 1315:23 2054:25]
  wire [3:0] _GEN_2239 = 7'h41 == cnt_layer ? 4'h0 : _GEN_2230; // @[control.scala 1315:23 2055:25]
  wire [7:0] _GEN_2240 = 7'h41 == cnt_layer ? 8'h0 : _GEN_2231; // @[control.scala 1315:23 2056:25]
  wire [7:0] _GEN_2241 = 7'h41 == cnt_layer ? 8'h0 : _GEN_2232; // @[control.scala 1315:23 2057:25]
  wire [31:0] _GEN_2242 = 7'h41 == cnt_layer ? 32'h3f800000 : _GEN_2233; // @[control.scala 1315:23 2058:25]
  wire [31:0] _GEN_2243 = 7'h41 == cnt_layer ? 32'h3f800000 : _GEN_2234; // @[control.scala 1315:23 2059:25]
  wire [7:0] _GEN_2244 = 7'h41 == cnt_layer ? 8'h0 : _GEN_2235; // @[control.scala 1315:23 2060:25]
  wire [31:0] _GEN_2245 = 7'h41 == cnt_layer ? 32'h22248000 : _GEN_2236; // @[control.scala 1315:23 2061:31]
  wire [31:0] _GEN_2246 = 7'h41 == cnt_layer ? 32'h22d18800 : _GEN_2237; // @[control.scala 1315:23 2062:31]
  wire [15:0] _GEN_2247 = 7'h40 == cnt_layer ? 16'h1 : _GEN_2238; // @[control.scala 1315:23 2043:25]
  wire [3:0] _GEN_2248 = 7'h40 == cnt_layer ? 4'h0 : _GEN_2239; // @[control.scala 1315:23 2044:25]
  wire [7:0] _GEN_2249 = 7'h40 == cnt_layer ? 8'h0 : _GEN_2240; // @[control.scala 1315:23 2045:25]
  wire [7:0] _GEN_2250 = 7'h40 == cnt_layer ? 8'h0 : _GEN_2241; // @[control.scala 1315:23 2046:25]
  wire [31:0] _GEN_2251 = 7'h40 == cnt_layer ? 32'h3f800000 : _GEN_2242; // @[control.scala 1315:23 2047:25]
  wire [31:0] _GEN_2252 = 7'h40 == cnt_layer ? 32'h3f800000 : _GEN_2243; // @[control.scala 1315:23 2048:25]
  wire [7:0] _GEN_2253 = 7'h40 == cnt_layer ? 8'h0 : _GEN_2244; // @[control.scala 1315:23 2049:25]
  wire [31:0] _GEN_2254 = 7'h40 == cnt_layer ? 32'h22200000 : _GEN_2245; // @[control.scala 1315:23 2050:31]
  wire [31:0] _GEN_2255 = 7'h40 == cnt_layer ? 32'h22d18000 : _GEN_2246; // @[control.scala 1315:23 2051:31]
  wire [15:0] _GEN_2256 = 7'h3f == cnt_layer ? 16'h1 : _GEN_2247; // @[control.scala 1315:23 2032:25]
  wire [3:0] _GEN_2257 = 7'h3f == cnt_layer ? 4'h0 : _GEN_2248; // @[control.scala 1315:23 2033:25]
  wire [7:0] _GEN_2258 = 7'h3f == cnt_layer ? 8'h0 : _GEN_2249; // @[control.scala 1315:23 2034:25]
  wire [7:0] _GEN_2259 = 7'h3f == cnt_layer ? 8'h0 : _GEN_2250; // @[control.scala 1315:23 2035:25]
  wire [31:0] _GEN_2260 = 7'h3f == cnt_layer ? 32'h3f800000 : _GEN_2251; // @[control.scala 1315:23 2036:25]
  wire [31:0] _GEN_2261 = 7'h3f == cnt_layer ? 32'h3f800000 : _GEN_2252; // @[control.scala 1315:23 2037:25]
  wire [7:0] _GEN_2262 = 7'h3f == cnt_layer ? 8'h0 : _GEN_2253; // @[control.scala 1315:23 2038:25]
  wire [31:0] _GEN_2263 = 7'h3f == cnt_layer ? 32'h221b8000 : _GEN_2254; // @[control.scala 1315:23 2039:31]
  wire [31:0] _GEN_2264 = 7'h3f == cnt_layer ? 32'h22d17800 : _GEN_2255; // @[control.scala 1315:23 2040:31]
  wire [15:0] _GEN_2265 = 7'h3e == cnt_layer ? 16'h1 : _GEN_2256; // @[control.scala 1315:23 2021:25]
  wire [3:0] _GEN_2266 = 7'h3e == cnt_layer ? 4'h0 : _GEN_2257; // @[control.scala 1315:23 2022:25]
  wire [7:0] _GEN_2267 = 7'h3e == cnt_layer ? 8'h0 : _GEN_2258; // @[control.scala 1315:23 2023:25]
  wire [7:0] _GEN_2268 = 7'h3e == cnt_layer ? 8'h0 : _GEN_2259; // @[control.scala 1315:23 2024:25]
  wire [31:0] _GEN_2269 = 7'h3e == cnt_layer ? 32'h3f800000 : _GEN_2260; // @[control.scala 1315:23 2025:25]
  wire [31:0] _GEN_2270 = 7'h3e == cnt_layer ? 32'h3f800000 : _GEN_2261; // @[control.scala 1315:23 2026:25]
  wire [7:0] _GEN_2271 = 7'h3e == cnt_layer ? 8'h0 : _GEN_2262; // @[control.scala 1315:23 2027:25]
  wire [31:0] _GEN_2272 = 7'h3e == cnt_layer ? 32'h22170000 : _GEN_2263; // @[control.scala 1315:23 2028:31]
  wire [31:0] _GEN_2273 = 7'h3e == cnt_layer ? 32'h22d17000 : _GEN_2264; // @[control.scala 1315:23 2029:31]
  wire [15:0] _GEN_2274 = 7'h3d == cnt_layer ? 16'h6544 : _GEN_2265; // @[control.scala 1315:23 2010:25]
  wire [3:0] _GEN_2275 = 7'h3d == cnt_layer ? 4'h8 : _GEN_2266; // @[control.scala 1315:23 2011:25]
  wire [7:0] _GEN_2276 = 7'h3d == cnt_layer ? 8'h6 : _GEN_2267; // @[control.scala 1315:23 2012:25]
  wire [7:0] _GEN_2277 = 7'h3d == cnt_layer ? 8'h40 : _GEN_2268; // @[control.scala 1315:23 2013:25]
  wire [31:0] _GEN_2278 = 7'h3d == cnt_layer ? 32'h3e184ea3 : _GEN_2269; // @[control.scala 1315:23 2014:25]
  wire [31:0] _GEN_2279 = 7'h3d == cnt_layer ? 32'h4153e89e : _GEN_2270; // @[control.scala 1315:23 2015:25]
  wire [7:0] _GEN_2280 = 7'h3d == cnt_layer ? 8'h4 : _GEN_2271; // @[control.scala 1315:23 2016:25]
  wire [31:0] _GEN_2281 = 7'h3d == cnt_layer ? 32'h22128000 : _GEN_2272; // @[control.scala 1315:23 2017:31]
  wire [31:0] _GEN_2282 = 7'h3d == cnt_layer ? 32'h22d16800 : _GEN_2273; // @[control.scala 1315:23 2018:31]
  wire [15:0] _GEN_2283 = 7'h3c == cnt_layer ? 16'h642b : _GEN_2274; // @[control.scala 1315:23 1999:25]
  wire [3:0] _GEN_2284 = 7'h3c == cnt_layer ? 4'h8 : _GEN_2275; // @[control.scala 1315:23 2000:25]
  wire [7:0] _GEN_2285 = 7'h3c == cnt_layer ? 8'h5 : _GEN_2276; // @[control.scala 1315:23 2001:25]
  wire [7:0] _GEN_2286 = 7'h3c == cnt_layer ? 8'h48 : _GEN_2277; // @[control.scala 1315:23 2002:25]
  wire [31:0] _GEN_2287 = 7'h3c == cnt_layer ? 32'h3dd6d44d : _GEN_2278; // @[control.scala 1315:23 2003:25]
  wire [31:0] _GEN_2288 = 7'h3c == cnt_layer ? 32'h41a9f3b9 : _GEN_2279; // @[control.scala 1315:23 2004:25]
  wire [7:0] _GEN_2289 = 7'h3c == cnt_layer ? 8'h6 : _GEN_2280; // @[control.scala 1315:23 2005:25]
  wire [31:0] _GEN_2290 = 7'h3c == cnt_layer ? 32'h220e0000 : _GEN_2281; // @[control.scala 1315:23 2006:31]
  wire [31:0] _GEN_2291 = 7'h3c == cnt_layer ? 32'h22d16000 : _GEN_2282; // @[control.scala 1315:23 2007:31]
  wire [15:0] _GEN_2292 = 7'h3b == cnt_layer ? 16'h4c2c : _GEN_2283; // @[control.scala 1315:23 1988:25]
  wire [3:0] _GEN_2293 = 7'h3b == cnt_layer ? 4'h7 : _GEN_2284; // @[control.scala 1315:23 1989:25]
  wire [7:0] _GEN_2294 = 7'h3b == cnt_layer ? 8'h3 : _GEN_2285; // @[control.scala 1315:23 1990:25]
  wire [7:0] _GEN_2295 = 7'h3b == cnt_layer ? 8'h52 : _GEN_2286; // @[control.scala 1315:23 1991:25]
  wire [31:0] _GEN_2296 = 7'h3b == cnt_layer ? 32'h3e21f651 : _GEN_2287; // @[control.scala 1315:23 1992:25]
  wire [31:0] _GEN_2297 = 7'h3b == cnt_layer ? 32'h4188e4c0 : _GEN_2288; // @[control.scala 1315:23 1993:25]
  wire [7:0] _GEN_2298 = 7'h3b == cnt_layer ? 8'h5 : _GEN_2289; // @[control.scala 1315:23 1994:25]
  wire [31:0] _GEN_2299 = 7'h3b == cnt_layer ? 32'h22098000 : _GEN_2290; // @[control.scala 1315:23 1995:31]
  wire [31:0] _GEN_2300 = 7'h3b == cnt_layer ? 32'h22d15800 : _GEN_2291; // @[control.scala 1315:23 1996:31]
  wire [15:0] _GEN_2301 = 7'h3a == cnt_layer ? 16'h43bc : _GEN_2292; // @[control.scala 1315:23 1975:25]
  wire [3:0] _GEN_2302 = 7'h3a == cnt_layer ? 4'h7 : _GEN_2293; // @[control.scala 1315:23 1976:25]
  wire [7:0] _GEN_2303 = 7'h3a == cnt_layer ? 8'h3 : _GEN_2294; // @[control.scala 1315:23 1977:25]
  wire [7:0] _GEN_2304 = 7'h3a == cnt_layer ? 8'h48 : _GEN_2295; // @[control.scala 1315:23 1978:25]
  wire [31:0] _GEN_2305 = 7'h3a == cnt_layer ? 32'h3e3d33de : _GEN_2296; // @[control.scala 1315:23 1979:25]
  wire [31:0] _GEN_2306 = 7'h3a == cnt_layer ? 32'h41415528 : _GEN_2297; // @[control.scala 1315:23 1980:25]
  wire [7:0] _GEN_2307 = 7'h3a == cnt_layer ? 8'h3 : _GEN_2298; // @[control.scala 1315:23 1981:25]
  wire [31:0] _GEN_2308 = 7'h3a == cnt_layer ? 32'h22050000 : _GEN_2299; // @[control.scala 1315:23 1982:31]
  wire [31:0] _GEN_2309 = 7'h3a == cnt_layer ? 32'h22d15000 : _GEN_2300; // @[control.scala 1315:23 1983:31]
  wire [15:0] _GEN_2310 = 7'h39 == cnt_layer ? 16'h1 : _GEN_2301; // @[control.scala 1315:23 1964:25]
  wire [3:0] _GEN_2311 = 7'h39 == cnt_layer ? 4'h0 : _GEN_2302; // @[control.scala 1315:23 1965:25]
  wire [7:0] _GEN_2312 = 7'h39 == cnt_layer ? 8'h0 : _GEN_2303; // @[control.scala 1315:23 1966:25]
  wire [7:0] _GEN_2313 = 7'h39 == cnt_layer ? 8'h0 : _GEN_2304; // @[control.scala 1315:23 1967:25]
  wire [31:0] _GEN_2314 = 7'h39 == cnt_layer ? 32'h3f800000 : _GEN_2305; // @[control.scala 1315:23 1968:25]
  wire [31:0] _GEN_2315 = 7'h39 == cnt_layer ? 32'h3f800000 : _GEN_2306; // @[control.scala 1315:23 1969:25]
  wire [7:0] _GEN_2316 = 7'h39 == cnt_layer ? 8'h0 : _GEN_2307; // @[control.scala 1315:23 1970:25]
  wire [31:0] _GEN_2317 = 7'h39 == cnt_layer ? 32'h22008000 : _GEN_2308; // @[control.scala 1315:23 1971:31]
  wire [31:0] _GEN_2318 = 7'h39 == cnt_layer ? 32'h22d14800 : _GEN_2309; // @[control.scala 1315:23 1972:31]
  wire [15:0] _GEN_2319 = 7'h38 == cnt_layer ? 16'h1 : _GEN_2310; // @[control.scala 1315:23 1953:25]
  wire [3:0] _GEN_2320 = 7'h38 == cnt_layer ? 4'h0 : _GEN_2311; // @[control.scala 1315:23 1954:25]
  wire [7:0] _GEN_2321 = 7'h38 == cnt_layer ? 8'h0 : _GEN_2312; // @[control.scala 1315:23 1955:25]
  wire [7:0] _GEN_2322 = 7'h38 == cnt_layer ? 8'h0 : _GEN_2313; // @[control.scala 1315:23 1956:25]
  wire [31:0] _GEN_2323 = 7'h38 == cnt_layer ? 32'h3f800000 : _GEN_2314; // @[control.scala 1315:23 1957:25]
  wire [31:0] _GEN_2324 = 7'h38 == cnt_layer ? 32'h3f800000 : _GEN_2315; // @[control.scala 1315:23 1958:25]
  wire [7:0] _GEN_2325 = 7'h38 == cnt_layer ? 8'h0 : _GEN_2316; // @[control.scala 1315:23 1959:25]
  wire [31:0] _GEN_2326 = 7'h38 == cnt_layer ? 32'h21fc0000 : _GEN_2317; // @[control.scala 1315:23 1960:31]
  wire [31:0] _GEN_2327 = 7'h38 == cnt_layer ? 32'h22d14000 : _GEN_2318; // @[control.scala 1315:23 1961:31]
  wire [15:0] _GEN_2328 = 7'h37 == cnt_layer ? 16'h1 : _GEN_2319; // @[control.scala 1315:23 1942:25]
  wire [3:0] _GEN_2329 = 7'h37 == cnt_layer ? 4'h0 : _GEN_2320; // @[control.scala 1315:23 1943:25]
  wire [7:0] _GEN_2330 = 7'h37 == cnt_layer ? 8'h0 : _GEN_2321; // @[control.scala 1315:23 1944:25]
  wire [7:0] _GEN_2331 = 7'h37 == cnt_layer ? 8'h0 : _GEN_2322; // @[control.scala 1315:23 1945:25]
  wire [31:0] _GEN_2332 = 7'h37 == cnt_layer ? 32'h3f800000 : _GEN_2323; // @[control.scala 1315:23 1946:25]
  wire [31:0] _GEN_2333 = 7'h37 == cnt_layer ? 32'h3f800000 : _GEN_2324; // @[control.scala 1315:23 1947:25]
  wire [7:0] _GEN_2334 = 7'h37 == cnt_layer ? 8'h0 : _GEN_2325; // @[control.scala 1315:23 1948:25]
  wire [31:0] _GEN_2335 = 7'h37 == cnt_layer ? 32'h21f78000 : _GEN_2326; // @[control.scala 1315:23 1949:31]
  wire [31:0] _GEN_2336 = 7'h37 == cnt_layer ? 32'h22d13800 : _GEN_2327; // @[control.scala 1315:23 1950:31]
  wire [15:0] _GEN_2337 = 7'h36 == cnt_layer ? 16'h1 : _GEN_2328; // @[control.scala 1315:23 1931:25]
  wire [3:0] _GEN_2338 = 7'h36 == cnt_layer ? 4'h0 : _GEN_2329; // @[control.scala 1315:23 1932:25]
  wire [7:0] _GEN_2339 = 7'h36 == cnt_layer ? 8'h0 : _GEN_2330; // @[control.scala 1315:23 1933:25]
  wire [7:0] _GEN_2340 = 7'h36 == cnt_layer ? 8'h0 : _GEN_2331; // @[control.scala 1315:23 1934:25]
  wire [31:0] _GEN_2341 = 7'h36 == cnt_layer ? 32'h3f800000 : _GEN_2332; // @[control.scala 1315:23 1935:25]
  wire [31:0] _GEN_2342 = 7'h36 == cnt_layer ? 32'h3f800000 : _GEN_2333; // @[control.scala 1315:23 1936:25]
  wire [7:0] _GEN_2343 = 7'h36 == cnt_layer ? 8'h0 : _GEN_2334; // @[control.scala 1315:23 1937:25]
  wire [31:0] _GEN_2344 = 7'h36 == cnt_layer ? 32'h21f30000 : _GEN_2335; // @[control.scala 1315:23 1938:31]
  wire [31:0] _GEN_2345 = 7'h36 == cnt_layer ? 32'h22d13000 : _GEN_2336; // @[control.scala 1315:23 1939:31]
  wire [15:0] _GEN_2346 = 7'h35 == cnt_layer ? 16'h451c : _GEN_2337; // @[control.scala 1315:23 1920:25]
  wire [3:0] _GEN_2347 = 7'h35 == cnt_layer ? 4'h7 : _GEN_2338; // @[control.scala 1315:23 1921:25]
  wire [7:0] _GEN_2348 = 7'h35 == cnt_layer ? 8'h4 : _GEN_2339; // @[control.scala 1315:23 1922:25]
  wire [7:0] _GEN_2349 = 7'h35 == cnt_layer ? 8'h3d : _GEN_2340; // @[control.scala 1315:23 1923:25]
  wire [31:0] _GEN_2350 = 7'h35 == cnt_layer ? 32'h3e262789 : _GEN_2341; // @[control.scala 1315:23 1924:25]
  wire [31:0] _GEN_2351 = 7'h35 == cnt_layer ? 32'h413950d9 : _GEN_2342; // @[control.scala 1315:23 1925:25]
  wire [7:0] _GEN_2352 = 7'h35 == cnt_layer ? 8'h3 : _GEN_2343; // @[control.scala 1315:23 1926:25]
  wire [31:0] _GEN_2353 = 7'h35 == cnt_layer ? 32'h21ee8000 : _GEN_2344; // @[control.scala 1315:23 1927:31]
  wire [31:0] _GEN_2354 = 7'h35 == cnt_layer ? 32'h22d12800 : _GEN_2345; // @[control.scala 1315:23 1928:31]
  wire [15:0] _GEN_2355 = 7'h34 == cnt_layer ? 16'h4b0f : _GEN_2346; // @[control.scala 1315:23 1909:25]
  wire [3:0] _GEN_2356 = 7'h34 == cnt_layer ? 4'h8 : _GEN_2347; // @[control.scala 1315:23 1910:25]
  wire [7:0] _GEN_2357 = 7'h34 == cnt_layer ? 8'h4 : _GEN_2348; // @[control.scala 1315:23 1911:25]
  wire [7:0] _GEN_2358 = 7'h34 == cnt_layer ? 8'h49 : _GEN_2349; // @[control.scala 1315:23 1912:25]
  wire [31:0] _GEN_2359 = 7'h34 == cnt_layer ? 32'h3e1c8b75 : _GEN_2350; // @[control.scala 1315:23 1913:25]
  wire [31:0] _GEN_2360 = 7'h34 == cnt_layer ? 32'h416dd3d5 : _GEN_2351; // @[control.scala 1315:23 1914:25]
  wire [7:0] _GEN_2361 = 7'h34 == cnt_layer ? 8'h4 : _GEN_2352; // @[control.scala 1315:23 1915:25]
  wire [31:0] _GEN_2362 = 7'h34 == cnt_layer ? 32'h21ea0000 : _GEN_2353; // @[control.scala 1315:23 1916:31]
  wire [31:0] _GEN_2363 = 7'h34 == cnt_layer ? 32'h22d12000 : _GEN_2354; // @[control.scala 1315:23 1917:31]
  wire [15:0] _GEN_2364 = 7'h33 == cnt_layer ? 16'h7b77 : _GEN_2355; // @[control.scala 1315:23 1898:25]
  wire [3:0] _GEN_2365 = 7'h33 == cnt_layer ? 4'h7 : _GEN_2356; // @[control.scala 1315:23 1899:25]
  wire [7:0] _GEN_2366 = 7'h33 == cnt_layer ? 8'h3 : _GEN_2357; // @[control.scala 1315:23 1900:25]
  wire [7:0] _GEN_2367 = 7'h33 == cnt_layer ? 8'h42 : _GEN_2358; // @[control.scala 1315:23 1901:25]
  wire [31:0] _GEN_2368 = 7'h33 == cnt_layer ? 32'h3e1ca663 : _GEN_2359; // @[control.scala 1315:23 1902:25]
  wire [31:0] _GEN_2369 = 7'h33 == cnt_layer ? 32'h41528e83 : _GEN_2360; // @[control.scala 1315:23 1903:25]
  wire [7:0] _GEN_2370 = 7'h33 == cnt_layer ? 8'h4 : _GEN_2361; // @[control.scala 1315:23 1904:25]
  wire [31:0] _GEN_2371 = 7'h33 == cnt_layer ? 32'h21e58000 : _GEN_2362; // @[control.scala 1315:23 1905:31]
  wire [31:0] _GEN_2372 = 7'h33 == cnt_layer ? 32'h22d11800 : _GEN_2363; // @[control.scala 1315:23 1906:31]
  wire [15:0] _GEN_2373 = 7'h32 == cnt_layer ? 16'h5f8a : _GEN_2364; // @[control.scala 1315:23 1886:24]
  wire [3:0] _GEN_2374 = 7'h32 == cnt_layer ? 4'h8 : _GEN_2365; // @[control.scala 1315:23 1887:24]
  wire [7:0] _GEN_2375 = 7'h32 == cnt_layer ? 8'h4 : _GEN_2366; // @[control.scala 1315:23 1888:19]
  wire [7:0] _GEN_2376 = 7'h32 == cnt_layer ? 8'h3b : _GEN_2367; // @[control.scala 1315:23 1889:20]
  wire [31:0] _GEN_2377 = 7'h32 == cnt_layer ? 32'h3e24718f : _GEN_2368; // @[control.scala 1315:23 1890:25]
  wire [31:0] _GEN_2378 = 7'h32 == cnt_layer ? 32'h4135f284 : _GEN_2369; // @[control.scala 1315:23 1891:25]
  wire [7:0] _GEN_2379 = 7'h32 == cnt_layer ? 8'h3 : _GEN_2370; // @[control.scala 1315:23 1892:20]
  wire [31:0] _GEN_2380 = 7'h32 == cnt_layer ? 32'h21e10000 : _GEN_2371; // @[control.scala 1315:23 1893:31]
  wire [31:0] _GEN_2381 = 7'h32 == cnt_layer ? 32'h22d11000 : _GEN_2372; // @[control.scala 1315:23 1894:31]
  wire [15:0] _GEN_2382 = 7'h31 == cnt_layer ? 16'h5a79 : _GEN_2373; // @[control.scala 1315:23 1875:24]
  wire [3:0] _GEN_2383 = 7'h31 == cnt_layer ? 4'h7 : _GEN_2374; // @[control.scala 1315:23 1876:24]
  wire [7:0] _GEN_2384 = 7'h31 == cnt_layer ? 8'h3 : _GEN_2375; // @[control.scala 1315:23 1877:19]
  wire [7:0] _GEN_2385 = 7'h31 == cnt_layer ? 8'h49 : _GEN_2376; // @[control.scala 1315:23 1878:20]
  wire [31:0] _GEN_2386 = 7'h31 == cnt_layer ? 32'h3e1baf4c : _GEN_2377; // @[control.scala 1315:23 1879:25]
  wire [31:0] _GEN_2387 = 7'h31 == cnt_layer ? 32'h417042cc : _GEN_2378; // @[control.scala 1315:23 1880:25]
  wire [7:0] _GEN_2388 = 7'h31 == cnt_layer ? 8'h4 : _GEN_2379; // @[control.scala 1315:23 1881:20]
  wire [31:0] _GEN_2389 = 7'h31 == cnt_layer ? 32'h21dc8000 : _GEN_2380; // @[control.scala 1315:23 1882:31]
  wire [31:0] _GEN_2390 = 7'h31 == cnt_layer ? 32'h22d10800 : _GEN_2381; // @[control.scala 1315:23 1883:31]
  wire [15:0] _GEN_2391 = 7'h30 == cnt_layer ? 16'h7a57 : _GEN_2382; // @[control.scala 1315:23 1862:24]
  wire [3:0] _GEN_2392 = 7'h30 == cnt_layer ? 4'h8 : _GEN_2383; // @[control.scala 1315:23 1863:24]
  wire [7:0] _GEN_2393 = 7'h30 == cnt_layer ? 8'h2 : _GEN_2384; // @[control.scala 1315:23 1864:19]
  wire [7:0] _GEN_2394 = 7'h30 == cnt_layer ? 8'h43 : _GEN_2385; // @[control.scala 1315:23 1865:20]
  wire [31:0] _GEN_2395 = 7'h30 == cnt_layer ? 32'h3e58089a : _GEN_2386; // @[control.scala 1315:23 1866:25]
  wire [31:0] _GEN_2396 = 7'h30 == cnt_layer ? 32'h411de732 : _GEN_2387; // @[control.scala 1315:23 1867:25]
  wire [7:0] _GEN_2397 = 7'h30 == cnt_layer ? 8'h3 : _GEN_2388; // @[control.scala 1315:23 1868:20]
  wire [31:0] _GEN_2398 = 7'h30 == cnt_layer ? 32'h21d80000 : _GEN_2389; // @[control.scala 1315:23 1869:31]
  wire [31:0] _GEN_2399 = 7'h30 == cnt_layer ? 32'h22d10000 : _GEN_2390; // @[control.scala 1315:23 1870:31]
  wire [15:0] _GEN_2400 = 7'h2f == cnt_layer ? 16'h1 : _GEN_2391; // @[control.scala 1315:23 1851:24]
  wire [3:0] _GEN_2401 = 7'h2f == cnt_layer ? 4'h0 : _GEN_2392; // @[control.scala 1315:23 1852:24]
  wire [7:0] _GEN_2402 = 7'h2f == cnt_layer ? 8'h0 : _GEN_2393; // @[control.scala 1315:23 1853:19]
  wire [7:0] _GEN_2403 = 7'h2f == cnt_layer ? 8'h0 : _GEN_2394; // @[control.scala 1315:23 1854:20]
  wire [31:0] _GEN_2404 = 7'h2f == cnt_layer ? 32'h3f800000 : _GEN_2395; // @[control.scala 1315:23 1855:25]
  wire [31:0] _GEN_2405 = 7'h2f == cnt_layer ? 32'h3f800000 : _GEN_2396; // @[control.scala 1315:23 1856:25]
  wire [7:0] _GEN_2406 = 7'h2f == cnt_layer ? 8'h0 : _GEN_2397; // @[control.scala 1315:23 1857:20]
  wire [31:0] _GEN_2407 = 7'h2f == cnt_layer ? 32'h21d38000 : _GEN_2398; // @[control.scala 1315:23 1858:31]
  wire [31:0] _GEN_2408 = 7'h2f == cnt_layer ? 32'h22d0f800 : _GEN_2399; // @[control.scala 1315:23 1859:31]
  wire [15:0] _GEN_2409 = 7'h2e == cnt_layer ? 16'h1 : _GEN_2400; // @[control.scala 1315:23 1840:24]
  wire [3:0] _GEN_2410 = 7'h2e == cnt_layer ? 4'h0 : _GEN_2401; // @[control.scala 1315:23 1841:24]
  wire [7:0] _GEN_2411 = 7'h2e == cnt_layer ? 8'h0 : _GEN_2402; // @[control.scala 1315:23 1842:19]
  wire [7:0] _GEN_2412 = 7'h2e == cnt_layer ? 8'h0 : _GEN_2403; // @[control.scala 1315:23 1843:20]
  wire [31:0] _GEN_2413 = 7'h2e == cnt_layer ? 32'h3f800000 : _GEN_2404; // @[control.scala 1315:23 1844:25]
  wire [31:0] _GEN_2414 = 7'h2e == cnt_layer ? 32'h3f800000 : _GEN_2405; // @[control.scala 1315:23 1845:25]
  wire [7:0] _GEN_2415 = 7'h2e == cnt_layer ? 8'h0 : _GEN_2406; // @[control.scala 1315:23 1846:20]
  wire [31:0] _GEN_2416 = 7'h2e == cnt_layer ? 32'h21cf0000 : _GEN_2407; // @[control.scala 1315:23 1847:31]
  wire [31:0] _GEN_2417 = 7'h2e == cnt_layer ? 32'h22d0f000 : _GEN_2408; // @[control.scala 1315:23 1848:31]
  wire [15:0] _GEN_2418 = 7'h2d == cnt_layer ? 16'h1 : _GEN_2409; // @[control.scala 1315:23 1829:24]
  wire [3:0] _GEN_2419 = 7'h2d == cnt_layer ? 4'h0 : _GEN_2410; // @[control.scala 1315:23 1830:24]
  wire [7:0] _GEN_2420 = 7'h2d == cnt_layer ? 8'h0 : _GEN_2411; // @[control.scala 1315:23 1831:19]
  wire [7:0] _GEN_2421 = 7'h2d == cnt_layer ? 8'h0 : _GEN_2412; // @[control.scala 1315:23 1832:20]
  wire [31:0] _GEN_2422 = 7'h2d == cnt_layer ? 32'h3f800000 : _GEN_2413; // @[control.scala 1315:23 1833:25]
  wire [31:0] _GEN_2423 = 7'h2d == cnt_layer ? 32'h3f800000 : _GEN_2414; // @[control.scala 1315:23 1834:25]
  wire [7:0] _GEN_2424 = 7'h2d == cnt_layer ? 8'h0 : _GEN_2415; // @[control.scala 1315:23 1835:20]
  wire [31:0] _GEN_2425 = 7'h2d == cnt_layer ? 32'h21ca8000 : _GEN_2416; // @[control.scala 1315:23 1836:31]
  wire [31:0] _GEN_2426 = 7'h2d == cnt_layer ? 32'h22d0e800 : _GEN_2417; // @[control.scala 1315:23 1837:31]
  wire [15:0] _GEN_2427 = 7'h2c == cnt_layer ? 16'h1 : _GEN_2418; // @[control.scala 1315:23 1818:24]
  wire [3:0] _GEN_2428 = 7'h2c == cnt_layer ? 4'h0 : _GEN_2419; // @[control.scala 1315:23 1819:24]
  wire [7:0] _GEN_2429 = 7'h2c == cnt_layer ? 8'h0 : _GEN_2420; // @[control.scala 1315:23 1820:19]
  wire [7:0] _GEN_2430 = 7'h2c == cnt_layer ? 8'h0 : _GEN_2421; // @[control.scala 1315:23 1821:20]
  wire [31:0] _GEN_2431 = 7'h2c == cnt_layer ? 32'h3f800000 : _GEN_2422; // @[control.scala 1315:23 1822:25]
  wire [31:0] _GEN_2432 = 7'h2c == cnt_layer ? 32'h3f800000 : _GEN_2423; // @[control.scala 1315:23 1823:25]
  wire [7:0] _GEN_2433 = 7'h2c == cnt_layer ? 8'h0 : _GEN_2424; // @[control.scala 1315:23 1824:20]
  wire [31:0] _GEN_2434 = 7'h2c == cnt_layer ? 32'h21c60000 : _GEN_2425; // @[control.scala 1315:23 1825:31]
  wire [31:0] _GEN_2435 = 7'h2c == cnt_layer ? 32'h22d0e000 : _GEN_2426; // @[control.scala 1315:23 1826:31]
  wire [15:0] _GEN_2436 = 7'h2b == cnt_layer ? 16'h5dc6 : _GEN_2427; // @[control.scala 1315:23 1807:24]
  wire [3:0] _GEN_2437 = 7'h2b == cnt_layer ? 4'h7 : _GEN_2428; // @[control.scala 1315:23 1808:24]
  wire [7:0] _GEN_2438 = 7'h2b == cnt_layer ? 8'h2 : _GEN_2429; // @[control.scala 1315:23 1809:19]
  wire [7:0] _GEN_2439 = 7'h2b == cnt_layer ? 8'h3e : _GEN_2430; // @[control.scala 1315:23 1810:20]
  wire [31:0] _GEN_2440 = 7'h2b == cnt_layer ? 32'h3e9db9c6 : _GEN_2431; // @[control.scala 1315:23 1811:25]
  wire [31:0] _GEN_2441 = 7'h2b == cnt_layer ? 32'h40c8f2a4 : _GEN_2432; // @[control.scala 1315:23 1812:25]
  wire [7:0] _GEN_2442 = 7'h2b == cnt_layer ? 8'h2 : _GEN_2433; // @[control.scala 1315:23 1813:20]
  wire [31:0] _GEN_2443 = 7'h2b == cnt_layer ? 32'h21c18000 : _GEN_2434; // @[control.scala 1315:23 1814:31]
  wire [31:0] _GEN_2444 = 7'h2b == cnt_layer ? 32'h22d0d800 : _GEN_2435; // @[control.scala 1315:23 1815:31]
  wire [15:0] _GEN_2445 = 7'h2a == cnt_layer ? 16'h41b5 : _GEN_2436; // @[control.scala 1315:23 1796:24]
  wire [3:0] _GEN_2446 = 7'h2a == cnt_layer ? 4'h7 : _GEN_2437; // @[control.scala 1315:23 1797:24]
  wire [7:0] _GEN_2447 = 7'h2a == cnt_layer ? 8'h2 : _GEN_2438; // @[control.scala 1315:23 1798:19]
  wire [7:0] _GEN_2448 = 7'h2a == cnt_layer ? 8'h39 : _GEN_2439; // @[control.scala 1315:23 1799:20]
  wire [31:0] _GEN_2449 = 7'h2a == cnt_layer ? 32'h3e76dc8e : _GEN_2440; // @[control.scala 1315:23 1800:25]
  wire [31:0] _GEN_2450 = 7'h2a == cnt_layer ? 32'h40eb7782 : _GEN_2441; // @[control.scala 1315:23 1801:25]
  wire [7:0] _GEN_2451 = 7'h2a == cnt_layer ? 8'h2 : _GEN_2442; // @[control.scala 1315:23 1802:20]
  wire [31:0] _GEN_2452 = 7'h2a == cnt_layer ? 32'h21bd0000 : _GEN_2443; // @[control.scala 1315:23 1803:31]
  wire [31:0] _GEN_2453 = 7'h2a == cnt_layer ? 32'h22d0d000 : _GEN_2444; // @[control.scala 1315:23 1804:31]
  wire [15:0] _GEN_2454 = 7'h29 == cnt_layer ? 16'h7a2a : _GEN_2445; // @[control.scala 1315:23 1785:24]
  wire [3:0] _GEN_2455 = 7'h29 == cnt_layer ? 4'h8 : _GEN_2446; // @[control.scala 1315:23 1786:24]
  wire [7:0] _GEN_2456 = 7'h29 == cnt_layer ? 8'h3 : _GEN_2447; // @[control.scala 1315:23 1787:19]
  wire [7:0] _GEN_2457 = 7'h29 == cnt_layer ? 8'h3a : _GEN_2448; // @[control.scala 1315:23 1788:20]
  wire [31:0] _GEN_2458 = 7'h29 == cnt_layer ? 32'h3e877345 : _GEN_2449; // @[control.scala 1315:23 1789:25]
  wire [31:0] _GEN_2459 = 7'h29 == cnt_layer ? 32'h40dc2a05 : _GEN_2450; // @[control.scala 1315:23 1790:25]
  wire [7:0] _GEN_2460 = 7'h29 == cnt_layer ? 8'h2 : _GEN_2451; // @[control.scala 1315:23 1791:20]
  wire [31:0] _GEN_2461 = 7'h29 == cnt_layer ? 32'h21b88000 : _GEN_2452; // @[control.scala 1315:23 1792:31]
  wire [31:0] _GEN_2462 = 7'h29 == cnt_layer ? 32'h22d0c800 : _GEN_2453; // @[control.scala 1315:23 1793:31]
  wire [15:0] _GEN_2463 = 7'h28 == cnt_layer ? 16'h4fcb : _GEN_2454; // @[control.scala 1315:23 1773:24]
  wire [3:0] _GEN_2464 = 7'h28 == cnt_layer ? 4'h8 : _GEN_2455; // @[control.scala 1315:23 1774:24]
  wire [7:0] _GEN_2465 = 7'h28 == cnt_layer ? 8'h3 : _GEN_2456; // @[control.scala 1315:23 1775:19]
  wire [7:0] _GEN_2466 = 7'h28 == cnt_layer ? 8'h40 : _GEN_2457; // @[control.scala 1315:23 1776:20]
  wire [31:0] _GEN_2467 = 7'h28 == cnt_layer ? 32'h3e2900ca : _GEN_2458; // @[control.scala 1315:23 1777:25]
  wire [31:0] _GEN_2468 = 7'h28 == cnt_layer ? 32'h413e64ce : _GEN_2459; // @[control.scala 1315:23 1778:25]
  wire [7:0] _GEN_2469 = 7'h28 == cnt_layer ? 8'h3 : _GEN_2460; // @[control.scala 1315:23 1779:20]
  wire [31:0] _GEN_2470 = 7'h28 == cnt_layer ? 32'h21b40000 : _GEN_2461; // @[control.scala 1315:23 1780:31]
  wire [31:0] _GEN_2471 = 7'h28 == cnt_layer ? 32'h22d0c000 : _GEN_2462; // @[control.scala 1315:23 1781:31]
  wire [15:0] _GEN_2472 = 7'h27 == cnt_layer ? 16'h4e9a : _GEN_2463; // @[control.scala 1315:23 1761:24]
  wire [3:0] _GEN_2473 = 7'h27 == cnt_layer ? 4'h7 : _GEN_2464; // @[control.scala 1315:23 1762:24]
  wire [7:0] _GEN_2474 = 7'h27 == cnt_layer ? 8'h1 : _GEN_2465; // @[control.scala 1315:23 1763:19]
  wire [7:0] _GEN_2475 = 7'h27 == cnt_layer ? 8'h3f : _GEN_2466; // @[control.scala 1315:23 1764:20]
  wire [31:0] _GEN_2476 = 7'h27 == cnt_layer ? 32'h3e2f0ff7 : _GEN_2467; // @[control.scala 1315:23 1765:25]
  wire [31:0] _GEN_2477 = 7'h27 == cnt_layer ? 32'h4134cc60 : _GEN_2468; // @[control.scala 1315:23 1766:25]
  wire [7:0] _GEN_2478 = 7'h27 == cnt_layer ? 8'h3 : _GEN_2469; // @[control.scala 1315:23 1767:20]
  wire [31:0] _GEN_2479 = 7'h27 == cnt_layer ? 32'h21af8000 : _GEN_2470; // @[control.scala 1315:23 1768:31]
  wire [31:0] _GEN_2480 = 7'h27 == cnt_layer ? 32'h22d0b800 : _GEN_2471; // @[control.scala 1315:23 1769:31]
  wire [15:0] _GEN_2481 = 7'h26 == cnt_layer ? 16'h1 : _GEN_2472; // @[control.scala 1315:23 1750:24]
  wire [3:0] _GEN_2482 = 7'h26 == cnt_layer ? 4'h0 : _GEN_2473; // @[control.scala 1315:23 1751:24]
  wire [7:0] _GEN_2483 = 7'h26 == cnt_layer ? 8'h0 : _GEN_2474; // @[control.scala 1315:23 1752:19]
  wire [7:0] _GEN_2484 = 7'h26 == cnt_layer ? 8'h0 : _GEN_2475; // @[control.scala 1315:23 1753:20]
  wire [31:0] _GEN_2485 = 7'h26 == cnt_layer ? 32'h3f800000 : _GEN_2476; // @[control.scala 1315:23 1754:25]
  wire [31:0] _GEN_2486 = 7'h26 == cnt_layer ? 32'h3f800000 : _GEN_2477; // @[control.scala 1315:23 1755:25]
  wire [7:0] _GEN_2487 = 7'h26 == cnt_layer ? 8'h0 : _GEN_2478; // @[control.scala 1315:23 1756:20]
  wire [31:0] _GEN_2488 = 7'h26 == cnt_layer ? 32'h21ab0000 : _GEN_2479; // @[control.scala 1315:23 1757:31]
  wire [31:0] _GEN_2489 = 7'h26 == cnt_layer ? 32'h22d0b000 : _GEN_2480; // @[control.scala 1315:23 1758:31]
  wire [15:0] _GEN_2490 = 7'h25 == cnt_layer ? 16'h1 : _GEN_2481; // @[control.scala 1315:23 1739:24]
  wire [3:0] _GEN_2491 = 7'h25 == cnt_layer ? 4'h0 : _GEN_2482; // @[control.scala 1315:23 1740:24]
  wire [7:0] _GEN_2492 = 7'h25 == cnt_layer ? 8'h0 : _GEN_2483; // @[control.scala 1315:23 1741:19]
  wire [7:0] _GEN_2493 = 7'h25 == cnt_layer ? 8'h0 : _GEN_2484; // @[control.scala 1315:23 1742:20]
  wire [31:0] _GEN_2494 = 7'h25 == cnt_layer ? 32'h3f800000 : _GEN_2485; // @[control.scala 1315:23 1743:25]
  wire [31:0] _GEN_2495 = 7'h25 == cnt_layer ? 32'h3f800000 : _GEN_2486; // @[control.scala 1315:23 1744:25]
  wire [7:0] _GEN_2496 = 7'h25 == cnt_layer ? 8'h0 : _GEN_2487; // @[control.scala 1315:23 1745:20]
  wire [31:0] _GEN_2497 = 7'h25 == cnt_layer ? 32'h21a68000 : _GEN_2488; // @[control.scala 1315:23 1746:31]
  wire [31:0] _GEN_2498 = 7'h25 == cnt_layer ? 32'h22d0a800 : _GEN_2489; // @[control.scala 1315:23 1747:31]
  wire [15:0] _GEN_2499 = 7'h24 == cnt_layer ? 16'h1 : _GEN_2490; // @[control.scala 1315:23 1728:24]
  wire [3:0] _GEN_2500 = 7'h24 == cnt_layer ? 4'h0 : _GEN_2491; // @[control.scala 1315:23 1729:24]
  wire [7:0] _GEN_2501 = 7'h24 == cnt_layer ? 8'h0 : _GEN_2492; // @[control.scala 1315:23 1730:19]
  wire [7:0] _GEN_2502 = 7'h24 == cnt_layer ? 8'h0 : _GEN_2493; // @[control.scala 1315:23 1731:20]
  wire [31:0] _GEN_2503 = 7'h24 == cnt_layer ? 32'h3f800000 : _GEN_2494; // @[control.scala 1315:23 1732:25]
  wire [31:0] _GEN_2504 = 7'h24 == cnt_layer ? 32'h3f800000 : _GEN_2495; // @[control.scala 1315:23 1733:25]
  wire [7:0] _GEN_2505 = 7'h24 == cnt_layer ? 8'h0 : _GEN_2496; // @[control.scala 1315:23 1734:20]
  wire [31:0] _GEN_2506 = 7'h24 == cnt_layer ? 32'h21a20000 : _GEN_2497; // @[control.scala 1315:23 1735:31]
  wire [31:0] _GEN_2507 = 7'h24 == cnt_layer ? 32'h22d0a000 : _GEN_2498; // @[control.scala 1315:23 1736:31]
  wire [15:0] _GEN_2508 = 7'h23 == cnt_layer ? 16'h1 : _GEN_2499; // @[control.scala 1315:23 1717:24]
  wire [3:0] _GEN_2509 = 7'h23 == cnt_layer ? 4'h0 : _GEN_2500; // @[control.scala 1315:23 1718:24]
  wire [7:0] _GEN_2510 = 7'h23 == cnt_layer ? 8'h0 : _GEN_2501; // @[control.scala 1315:23 1719:19]
  wire [7:0] _GEN_2511 = 7'h23 == cnt_layer ? 8'h0 : _GEN_2502; // @[control.scala 1315:23 1720:20]
  wire [31:0] _GEN_2512 = 7'h23 == cnt_layer ? 32'h3f800000 : _GEN_2503; // @[control.scala 1315:23 1721:25]
  wire [31:0] _GEN_2513 = 7'h23 == cnt_layer ? 32'h3f800000 : _GEN_2504; // @[control.scala 1315:23 1722:25]
  wire [7:0] _GEN_2514 = 7'h23 == cnt_layer ? 8'h0 : _GEN_2505; // @[control.scala 1315:23 1723:20]
  wire [31:0] _GEN_2515 = 7'h23 == cnt_layer ? 32'h219d8000 : _GEN_2506; // @[control.scala 1315:23 1724:31]
  wire [31:0] _GEN_2516 = 7'h23 == cnt_layer ? 32'h22d09800 : _GEN_2507; // @[control.scala 1315:23 1725:31]
  wire [15:0] _GEN_2517 = 7'h22 == cnt_layer ? 16'h1 : _GEN_2508; // @[control.scala 1315:23 1706:24]
  wire [3:0] _GEN_2518 = 7'h22 == cnt_layer ? 4'h0 : _GEN_2509; // @[control.scala 1315:23 1707:24]
  wire [7:0] _GEN_2519 = 7'h22 == cnt_layer ? 8'h0 : _GEN_2510; // @[control.scala 1315:23 1708:19]
  wire [7:0] _GEN_2520 = 7'h22 == cnt_layer ? 8'h0 : _GEN_2511; // @[control.scala 1315:23 1709:20]
  wire [31:0] _GEN_2521 = 7'h22 == cnt_layer ? 32'h3f800000 : _GEN_2512; // @[control.scala 1315:23 1710:25]
  wire [31:0] _GEN_2522 = 7'h22 == cnt_layer ? 32'h3f800000 : _GEN_2513; // @[control.scala 1315:23 1711:25]
  wire [7:0] _GEN_2523 = 7'h22 == cnt_layer ? 8'h0 : _GEN_2514; // @[control.scala 1315:23 1712:20]
  wire [31:0] _GEN_2524 = 7'h22 == cnt_layer ? 32'h21990000 : _GEN_2515; // @[control.scala 1315:23 1713:31]
  wire [31:0] _GEN_2525 = 7'h22 == cnt_layer ? 32'h22d09000 : _GEN_2516; // @[control.scala 1315:23 1714:31]
  wire [15:0] _GEN_2526 = 7'h21 == cnt_layer ? 16'h1 : _GEN_2517; // @[control.scala 1315:23 1695:24]
  wire [3:0] _GEN_2527 = 7'h21 == cnt_layer ? 4'h0 : _GEN_2518; // @[control.scala 1315:23 1696:24]
  wire [7:0] _GEN_2528 = 7'h21 == cnt_layer ? 8'h0 : _GEN_2519; // @[control.scala 1315:23 1697:19]
  wire [7:0] _GEN_2529 = 7'h21 == cnt_layer ? 8'h0 : _GEN_2520; // @[control.scala 1315:23 1698:20]
  wire [31:0] _GEN_2530 = 7'h21 == cnt_layer ? 32'h3f800000 : _GEN_2521; // @[control.scala 1315:23 1699:25]
  wire [31:0] _GEN_2531 = 7'h21 == cnt_layer ? 32'h3f800000 : _GEN_2522; // @[control.scala 1315:23 1700:25]
  wire [7:0] _GEN_2532 = 7'h21 == cnt_layer ? 8'h0 : _GEN_2523; // @[control.scala 1315:23 1701:20]
  wire [31:0] _GEN_2533 = 7'h21 == cnt_layer ? 32'h21948000 : _GEN_2524; // @[control.scala 1315:23 1702:31]
  wire [31:0] _GEN_2534 = 7'h21 == cnt_layer ? 32'h22d08800 : _GEN_2525; // @[control.scala 1315:23 1703:31]
  wire [15:0] _GEN_2535 = 7'h20 == cnt_layer ? 16'h1 : _GEN_2526; // @[control.scala 1315:23 1684:24]
  wire [3:0] _GEN_2536 = 7'h20 == cnt_layer ? 4'h0 : _GEN_2527; // @[control.scala 1315:23 1685:24]
  wire [7:0] _GEN_2537 = 7'h20 == cnt_layer ? 8'h0 : _GEN_2528; // @[control.scala 1315:23 1686:19]
  wire [7:0] _GEN_2538 = 7'h20 == cnt_layer ? 8'h0 : _GEN_2529; // @[control.scala 1315:23 1687:20]
  wire [31:0] _GEN_2539 = 7'h20 == cnt_layer ? 32'h3f800000 : _GEN_2530; // @[control.scala 1315:23 1688:25]
  wire [31:0] _GEN_2540 = 7'h20 == cnt_layer ? 32'h3f800000 : _GEN_2531; // @[control.scala 1315:23 1689:25]
  wire [7:0] _GEN_2541 = 7'h20 == cnt_layer ? 8'h0 : _GEN_2532; // @[control.scala 1315:23 1690:20]
  wire [31:0] _GEN_2542 = 7'h20 == cnt_layer ? 32'h21900000 : _GEN_2533; // @[control.scala 1315:23 1691:31]
  wire [31:0] _GEN_2543 = 7'h20 == cnt_layer ? 32'h22d08000 : _GEN_2534; // @[control.scala 1315:23 1692:31]
  wire [15:0] _GEN_2544 = 7'h1f == cnt_layer ? 16'h1 : _GEN_2535; // @[control.scala 1315:23 1673:24]
  wire [3:0] _GEN_2545 = 7'h1f == cnt_layer ? 4'h0 : _GEN_2536; // @[control.scala 1315:23 1674:24]
  wire [7:0] _GEN_2546 = 7'h1f == cnt_layer ? 8'h0 : _GEN_2537; // @[control.scala 1315:23 1675:19]
  wire [7:0] _GEN_2547 = 7'h1f == cnt_layer ? 8'h0 : _GEN_2538; // @[control.scala 1315:23 1676:20]
  wire [31:0] _GEN_2548 = 7'h1f == cnt_layer ? 32'h3f800000 : _GEN_2539; // @[control.scala 1315:23 1677:25]
  wire [31:0] _GEN_2549 = 7'h1f == cnt_layer ? 32'h3f800000 : _GEN_2540; // @[control.scala 1315:23 1678:25]
  wire [7:0] _GEN_2550 = 7'h1f == cnt_layer ? 8'h0 : _GEN_2541; // @[control.scala 1315:23 1679:20]
  wire [31:0] _GEN_2551 = 7'h1f == cnt_layer ? 32'h218b8000 : _GEN_2542; // @[control.scala 1315:23 1680:31]
  wire [31:0] _GEN_2552 = 7'h1f == cnt_layer ? 32'h22d07800 : _GEN_2543; // @[control.scala 1315:23 1681:31]
  wire [15:0] _GEN_2553 = 7'h1e == cnt_layer ? 16'h5f2d : _GEN_2544; // @[control.scala 1315:23 1662:24]
  wire [3:0] _GEN_2554 = 7'h1e == cnt_layer ? 4'h7 : _GEN_2545; // @[control.scala 1315:23 1663:24]
  wire [7:0] _GEN_2555 = 7'h1e == cnt_layer ? 8'h3 : _GEN_2546; // @[control.scala 1315:23 1664:19]
  wire [7:0] _GEN_2556 = 7'h1e == cnt_layer ? 8'h32 : _GEN_2547; // @[control.scala 1315:23 1665:20]
  wire [31:0] _GEN_2557 = 7'h1e == cnt_layer ? 32'h3eabd6d9 : _GEN_2548; // @[control.scala 1315:23 1666:25]
  wire [31:0] _GEN_2558 = 7'h1e == cnt_layer ? 32'h409ac75f : _GEN_2549; // @[control.scala 1315:23 1667:25]
  wire [7:0] _GEN_2559 = 7'h1e == cnt_layer ? 8'h1 : _GEN_2550; // @[control.scala 1315:23 1668:20]
  wire [31:0] _GEN_2560 = 7'h1e == cnt_layer ? 32'h21870000 : _GEN_2551; // @[control.scala 1315:23 1669:31]
  wire [31:0] _GEN_2561 = 7'h1e == cnt_layer ? 32'h22d07000 : _GEN_2552; // @[control.scala 1315:23 1670:31]
  wire [15:0] _GEN_2562 = 7'h1d == cnt_layer ? 16'h543f : _GEN_2553; // @[control.scala 1315:23 1651:24]
  wire [3:0] _GEN_2563 = 7'h1d == cnt_layer ? 4'h8 : _GEN_2554; // @[control.scala 1315:23 1652:24]
  wire [7:0] _GEN_2564 = 7'h1d == cnt_layer ? 8'h4 : _GEN_2555; // @[control.scala 1315:23 1653:19]
  wire [7:0] _GEN_2565 = 7'h1d == cnt_layer ? 8'h34 : _GEN_2556; // @[control.scala 1315:23 1654:20]
  wire [31:0] _GEN_2566 = 7'h1d == cnt_layer ? 32'h3e2dff7e : _GEN_2557; // @[control.scala 1315:23 1655:25]
  wire [31:0] _GEN_2567 = 7'h1d == cnt_layer ? 32'h411c9ff6 : _GEN_2558; // @[control.scala 1315:23 1656:25]
  wire [7:0] _GEN_2568 = 7'h1d == cnt_layer ? 8'h3 : _GEN_2559; // @[control.scala 1315:23 1657:20]
  wire [31:0] _GEN_2569 = 7'h1d == cnt_layer ? 32'h21828000 : _GEN_2560; // @[control.scala 1315:23 1658:31]
  wire [31:0] _GEN_2570 = 7'h1d == cnt_layer ? 32'h22d06800 : _GEN_2561; // @[control.scala 1315:23 1659:31]
  wire [15:0] _GEN_2571 = 7'h1c == cnt_layer ? 16'h6c21 : _GEN_2562; // @[control.scala 1315:23 1640:24]
  wire [3:0] _GEN_2572 = 7'h1c == cnt_layer ? 4'h8 : _GEN_2563; // @[control.scala 1315:23 1641:24]
  wire [7:0] _GEN_2573 = 7'h1c == cnt_layer ? 8'h4 : _GEN_2564; // @[control.scala 1315:23 1642:19]
  wire [7:0] _GEN_2574 = 7'h1c == cnt_layer ? 8'h41 : _GEN_2565; // @[control.scala 1315:23 1643:20]
  wire [31:0] _GEN_2575 = 7'h1c == cnt_layer ? 32'h3e1744c8 : _GEN_2566; // @[control.scala 1315:23 1644:25]
  wire [31:0] _GEN_2576 = 7'h1c == cnt_layer ? 32'h41584614 : _GEN_2567; // @[control.scala 1315:23 1645:25]
  wire [7:0] _GEN_2577 = 7'h1c == cnt_layer ? 8'h4 : _GEN_2568; // @[control.scala 1315:23 1646:20]
  wire [31:0] _GEN_2578 = 7'h1c == cnt_layer ? 32'h217e0000 : _GEN_2569; // @[control.scala 1315:23 1647:31]
  wire [31:0] _GEN_2579 = 7'h1c == cnt_layer ? 32'h22d06000 : _GEN_2570; // @[control.scala 1315:23 1648:31]
  wire [15:0] _GEN_2580 = 7'h1b == cnt_layer ? 16'h5aa2 : _GEN_2571; // @[control.scala 1315:23 1629:24]
  wire [3:0] _GEN_2581 = 7'h1b == cnt_layer ? 4'h7 : _GEN_2572; // @[control.scala 1315:23 1630:24]
  wire [7:0] _GEN_2582 = 7'h1b == cnt_layer ? 8'h3 : _GEN_2573; // @[control.scala 1315:23 1631:19]
  wire [7:0] _GEN_2583 = 7'h1b == cnt_layer ? 8'h45 : _GEN_2574; // @[control.scala 1315:23 1632:20]
  wire [31:0] _GEN_2584 = 7'h1b == cnt_layer ? 32'h3e27474e : _GEN_2575; // @[control.scala 1315:23 1633:25]
  wire [31:0] _GEN_2585 = 7'h1b == cnt_layer ? 32'h41514282 : _GEN_2576; // @[control.scala 1315:23 1634:25]
  wire [7:0] _GEN_2586 = 7'h1b == cnt_layer ? 8'h4 : _GEN_2577; // @[control.scala 1315:23 1635:20]
  wire [31:0] _GEN_2587 = 7'h1b == cnt_layer ? 32'h21798000 : _GEN_2578; // @[control.scala 1315:23 1636:31]
  wire [31:0] _GEN_2588 = 7'h1b == cnt_layer ? 32'h22d05800 : _GEN_2579; // @[control.scala 1315:23 1637:31]
  wire [15:0] _GEN_2589 = 7'h1a == cnt_layer ? 16'h66a0 : _GEN_2580; // @[control.scala 1315:23 1618:24]
  wire [3:0] _GEN_2590 = 7'h1a == cnt_layer ? 4'h7 : _GEN_2581; // @[control.scala 1315:23 1619:24]
  wire [7:0] _GEN_2591 = 7'h1a == cnt_layer ? 8'h4 : _GEN_2582; // @[control.scala 1315:23 1620:19]
  wire [7:0] _GEN_2592 = 7'h1a == cnt_layer ? 8'h49 : _GEN_2583; // @[control.scala 1315:23 1621:20]
  wire [31:0] _GEN_2593 = 7'h1a == cnt_layer ? 32'h3e3d9e99 : _GEN_2584; // @[control.scala 1315:23 1622:25]
  wire [31:0] _GEN_2594 = 7'h1a == cnt_layer ? 32'h4144788f : _GEN_2585; // @[control.scala 1315:23 1623:25]
  wire [7:0] _GEN_2595 = 7'h1a == cnt_layer ? 8'h3 : _GEN_2586; // @[control.scala 1315:23 1624:20]
  wire [31:0] _GEN_2596 = 7'h1a == cnt_layer ? 32'h21750000 : _GEN_2587; // @[control.scala 1315:23 1625:31]
  wire [31:0] _GEN_2597 = 7'h1a == cnt_layer ? 32'h22d05000 : _GEN_2588; // @[control.scala 1315:23 1626:31]
  wire [15:0] _GEN_2598 = 7'h19 == cnt_layer ? 16'h55c7 : _GEN_2589; // @[control.scala 1315:23 1606:24]
  wire [3:0] _GEN_2599 = 7'h19 == cnt_layer ? 4'h8 : _GEN_2590; // @[control.scala 1315:23 1607:24]
  wire [7:0] _GEN_2600 = 7'h19 == cnt_layer ? 8'h3 : _GEN_2591; // @[control.scala 1315:23 1608:19]
  wire [7:0] _GEN_2601 = 7'h19 == cnt_layer ? 8'h53 : _GEN_2592; // @[control.scala 1315:23 1609:20]
  wire [31:0] _GEN_2602 = 7'h19 == cnt_layer ? 32'h3e4825a3 : _GEN_2593; // @[control.scala 1315:23 1610:25]
  wire [31:0] _GEN_2603 = 7'h19 == cnt_layer ? 32'h416423c6 : _GEN_2594; // @[control.scala 1315:23 1611:25]
  wire [7:0] _GEN_2604 = 7'h19 == cnt_layer ? 8'h4 : _GEN_2595; // @[control.scala 1315:23 1612:20]
  wire [31:0] _GEN_2605 = 7'h19 == cnt_layer ? 32'h21708000 : _GEN_2596; // @[control.scala 1315:23 1613:31]
  wire [31:0] _GEN_2606 = 7'h19 == cnt_layer ? 32'h22d04800 : _GEN_2597; // @[control.scala 1315:23 1614:31]
  wire [15:0] _GEN_2607 = 7'h18 == cnt_layer ? 16'h5fe8 : _GEN_2598; // @[control.scala 1315:23 1594:24]
  wire [3:0] _GEN_2608 = 7'h18 == cnt_layer ? 4'h8 : _GEN_2599; // @[control.scala 1315:23 1595:24]
  wire [7:0] _GEN_2609 = 7'h18 == cnt_layer ? 8'h3 : _GEN_2600; // @[control.scala 1315:23 1596:19]
  wire [7:0] _GEN_2610 = 7'h18 == cnt_layer ? 8'h3e : _GEN_2601; // @[control.scala 1315:23 1597:20]
  wire [31:0] _GEN_2611 = 7'h18 == cnt_layer ? 32'h3e3e0a9b : _GEN_2602; // @[control.scala 1315:23 1598:25]
  wire [31:0] _GEN_2612 = 7'h18 == cnt_layer ? 32'h4123b903 : _GEN_2603; // @[control.scala 1315:23 1599:25]
  wire [7:0] _GEN_2613 = 7'h18 == cnt_layer ? 8'h3 : _GEN_2604; // @[control.scala 1315:23 1600:20]
  wire [31:0] _GEN_2614 = 7'h18 == cnt_layer ? 32'h216c0000 : _GEN_2605; // @[control.scala 1315:23 1601:31]
  wire [31:0] _GEN_2615 = 7'h18 == cnt_layer ? 32'h22d04000 : _GEN_2606; // @[control.scala 1315:23 1602:31]
  wire [15:0] _GEN_2616 = 7'h17 == cnt_layer ? 16'h1 : _GEN_2607; // @[control.scala 1315:23 1583:24]
  wire [3:0] _GEN_2617 = 7'h17 == cnt_layer ? 4'h0 : _GEN_2608; // @[control.scala 1315:23 1584:24]
  wire [7:0] _GEN_2618 = 7'h17 == cnt_layer ? 8'h0 : _GEN_2609; // @[control.scala 1315:23 1585:19]
  wire [7:0] _GEN_2619 = 7'h17 == cnt_layer ? 8'h0 : _GEN_2610; // @[control.scala 1315:23 1586:20]
  wire [31:0] _GEN_2620 = 7'h17 == cnt_layer ? 32'h3f800000 : _GEN_2611; // @[control.scala 1315:23 1587:25]
  wire [31:0] _GEN_2621 = 7'h17 == cnt_layer ? 32'h3f800000 : _GEN_2612; // @[control.scala 1315:23 1588:25]
  wire [7:0] _GEN_2622 = 7'h17 == cnt_layer ? 8'h0 : _GEN_2613; // @[control.scala 1315:23 1589:20]
  wire [31:0] _GEN_2623 = 7'h17 == cnt_layer ? 32'h21678000 : _GEN_2614; // @[control.scala 1315:23 1590:31]
  wire [31:0] _GEN_2624 = 7'h17 == cnt_layer ? 32'h22d03800 : _GEN_2615; // @[control.scala 1315:23 1591:31]
  wire [15:0] _GEN_2625 = 7'h16 == cnt_layer ? 16'h1 : _GEN_2616; // @[control.scala 1315:23 1572:24]
  wire [3:0] _GEN_2626 = 7'h16 == cnt_layer ? 4'h0 : _GEN_2617; // @[control.scala 1315:23 1573:24]
  wire [7:0] _GEN_2627 = 7'h16 == cnt_layer ? 8'h0 : _GEN_2618; // @[control.scala 1315:23 1574:19]
  wire [7:0] _GEN_2628 = 7'h16 == cnt_layer ? 8'h0 : _GEN_2619; // @[control.scala 1315:23 1575:20]
  wire [31:0] _GEN_2629 = 7'h16 == cnt_layer ? 32'h3f800000 : _GEN_2620; // @[control.scala 1315:23 1576:25]
  wire [31:0] _GEN_2630 = 7'h16 == cnt_layer ? 32'h3f800000 : _GEN_2621; // @[control.scala 1315:23 1577:25]
  wire [7:0] _GEN_2631 = 7'h16 == cnt_layer ? 8'h0 : _GEN_2622; // @[control.scala 1315:23 1578:20]
  wire [31:0] _GEN_2632 = 7'h16 == cnt_layer ? 32'h21630000 : _GEN_2623; // @[control.scala 1315:23 1579:31]
  wire [31:0] _GEN_2633 = 7'h16 == cnt_layer ? 32'h22d03000 : _GEN_2624; // @[control.scala 1315:23 1580:31]
  wire [15:0] _GEN_2634 = 7'h15 == cnt_layer ? 16'h1 : _GEN_2625; // @[control.scala 1315:23 1561:24]
  wire [3:0] _GEN_2635 = 7'h15 == cnt_layer ? 4'h0 : _GEN_2626; // @[control.scala 1315:23 1562:24]
  wire [7:0] _GEN_2636 = 7'h15 == cnt_layer ? 8'h0 : _GEN_2627; // @[control.scala 1315:23 1563:19]
  wire [7:0] _GEN_2637 = 7'h15 == cnt_layer ? 8'h0 : _GEN_2628; // @[control.scala 1315:23 1564:20]
  wire [31:0] _GEN_2638 = 7'h15 == cnt_layer ? 32'h3f800000 : _GEN_2629; // @[control.scala 1315:23 1565:25]
  wire [31:0] _GEN_2639 = 7'h15 == cnt_layer ? 32'h3f800000 : _GEN_2630; // @[control.scala 1315:23 1566:25]
  wire [7:0] _GEN_2640 = 7'h15 == cnt_layer ? 8'h0 : _GEN_2631; // @[control.scala 1315:23 1567:20]
  wire [31:0] _GEN_2641 = 7'h15 == cnt_layer ? 32'h215e8000 : _GEN_2632; // @[control.scala 1315:23 1568:31]
  wire [31:0] _GEN_2642 = 7'h15 == cnt_layer ? 32'h22d02800 : _GEN_2633; // @[control.scala 1315:23 1569:31]
  wire [15:0] _GEN_2643 = 7'h14 == cnt_layer ? 16'h1 : _GEN_2634; // @[control.scala 1315:23 1550:24]
  wire [3:0] _GEN_2644 = 7'h14 == cnt_layer ? 4'h0 : _GEN_2635; // @[control.scala 1315:23 1551:24]
  wire [7:0] _GEN_2645 = 7'h14 == cnt_layer ? 8'h0 : _GEN_2636; // @[control.scala 1315:23 1552:19]
  wire [7:0] _GEN_2646 = 7'h14 == cnt_layer ? 8'h0 : _GEN_2637; // @[control.scala 1315:23 1553:20]
  wire [31:0] _GEN_2647 = 7'h14 == cnt_layer ? 32'h3f800000 : _GEN_2638; // @[control.scala 1315:23 1554:25]
  wire [31:0] _GEN_2648 = 7'h14 == cnt_layer ? 32'h3f800000 : _GEN_2639; // @[control.scala 1315:23 1555:25]
  wire [7:0] _GEN_2649 = 7'h14 == cnt_layer ? 8'h0 : _GEN_2640; // @[control.scala 1315:23 1556:20]
  wire [31:0] _GEN_2650 = 7'h14 == cnt_layer ? 32'h215a0000 : _GEN_2641; // @[control.scala 1315:23 1557:31]
  wire [31:0] _GEN_2651 = 7'h14 == cnt_layer ? 32'h22d02000 : _GEN_2642; // @[control.scala 1315:23 1558:31]
  wire [15:0] _GEN_2652 = 7'h13 == cnt_layer ? 16'h1 : _GEN_2643; // @[control.scala 1315:23 1539:24]
  wire [3:0] _GEN_2653 = 7'h13 == cnt_layer ? 4'h0 : _GEN_2644; // @[control.scala 1315:23 1540:24]
  wire [7:0] _GEN_2654 = 7'h13 == cnt_layer ? 8'h0 : _GEN_2645; // @[control.scala 1315:23 1541:19]
  wire [7:0] _GEN_2655 = 7'h13 == cnt_layer ? 8'h0 : _GEN_2646; // @[control.scala 1315:23 1542:20]
  wire [31:0] _GEN_2656 = 7'h13 == cnt_layer ? 32'h3f800000 : _GEN_2647; // @[control.scala 1315:23 1543:25]
  wire [31:0] _GEN_2657 = 7'h13 == cnt_layer ? 32'h3f800000 : _GEN_2648; // @[control.scala 1315:23 1544:25]
  wire [7:0] _GEN_2658 = 7'h13 == cnt_layer ? 8'h0 : _GEN_2649; // @[control.scala 1315:23 1545:20]
  wire [31:0] _GEN_2659 = 7'h13 == cnt_layer ? 32'h21558000 : _GEN_2650; // @[control.scala 1315:23 1546:31]
  wire [31:0] _GEN_2660 = 7'h13 == cnt_layer ? 32'h22d01800 : _GEN_2651; // @[control.scala 1315:23 1547:31]
  wire [15:0] _GEN_2661 = 7'h12 == cnt_layer ? 16'h1 : _GEN_2652; // @[control.scala 1315:23 1528:24]
  wire [3:0] _GEN_2662 = 7'h12 == cnt_layer ? 4'h0 : _GEN_2653; // @[control.scala 1315:23 1529:24]
  wire [7:0] _GEN_2663 = 7'h12 == cnt_layer ? 8'h0 : _GEN_2654; // @[control.scala 1315:23 1530:19]
  wire [7:0] _GEN_2664 = 7'h12 == cnt_layer ? 8'h0 : _GEN_2655; // @[control.scala 1315:23 1531:20]
  wire [31:0] _GEN_2665 = 7'h12 == cnt_layer ? 32'h3f800000 : _GEN_2656; // @[control.scala 1315:23 1532:25]
  wire [31:0] _GEN_2666 = 7'h12 == cnt_layer ? 32'h3f800000 : _GEN_2657; // @[control.scala 1315:23 1533:25]
  wire [7:0] _GEN_2667 = 7'h12 == cnt_layer ? 8'h0 : _GEN_2658; // @[control.scala 1315:23 1534:20]
  wire [31:0] _GEN_2668 = 7'h12 == cnt_layer ? 32'h21510000 : _GEN_2659; // @[control.scala 1315:23 1535:31]
  wire [31:0] _GEN_2669 = 7'h12 == cnt_layer ? 32'h22d01000 : _GEN_2660; // @[control.scala 1315:23 1536:31]
  wire [15:0] _GEN_2670 = 7'h11 == cnt_layer ? 16'h1 : _GEN_2661; // @[control.scala 1315:23 1517:24]
  wire [3:0] _GEN_2671 = 7'h11 == cnt_layer ? 4'h0 : _GEN_2662; // @[control.scala 1315:23 1518:24]
  wire [7:0] _GEN_2672 = 7'h11 == cnt_layer ? 8'h0 : _GEN_2663; // @[control.scala 1315:23 1519:19]
  wire [7:0] _GEN_2673 = 7'h11 == cnt_layer ? 8'h0 : _GEN_2664; // @[control.scala 1315:23 1520:20]
  wire [31:0] _GEN_2674 = 7'h11 == cnt_layer ? 32'h3f800000 : _GEN_2665; // @[control.scala 1315:23 1521:25]
  wire [31:0] _GEN_2675 = 7'h11 == cnt_layer ? 32'h3f800000 : _GEN_2666; // @[control.scala 1315:23 1522:25]
  wire [7:0] _GEN_2676 = 7'h11 == cnt_layer ? 8'h0 : _GEN_2667; // @[control.scala 1315:23 1523:20]
  wire [31:0] _GEN_2677 = 7'h11 == cnt_layer ? 32'h214c8000 : _GEN_2668; // @[control.scala 1315:23 1524:31]
  wire [31:0] _GEN_2678 = 7'h11 == cnt_layer ? 32'h22d00800 : _GEN_2669; // @[control.scala 1315:23 1525:31]
  wire [15:0] _GEN_2679 = 7'h10 == cnt_layer ? 16'h1 : _GEN_2670; // @[control.scala 1315:23 1506:24]
  wire [3:0] _GEN_2680 = 7'h10 == cnt_layer ? 4'h0 : _GEN_2671; // @[control.scala 1315:23 1507:24]
  wire [7:0] _GEN_2681 = 7'h10 == cnt_layer ? 8'h0 : _GEN_2672; // @[control.scala 1315:23 1508:19]
  wire [7:0] _GEN_2682 = 7'h10 == cnt_layer ? 8'h0 : _GEN_2673; // @[control.scala 1315:23 1509:20]
  wire [31:0] _GEN_2683 = 7'h10 == cnt_layer ? 32'h3f800000 : _GEN_2674; // @[control.scala 1315:23 1510:25]
  wire [31:0] _GEN_2684 = 7'h10 == cnt_layer ? 32'h3f800000 : _GEN_2675; // @[control.scala 1315:23 1511:25]
  wire [7:0] _GEN_2685 = 7'h10 == cnt_layer ? 8'h0 : _GEN_2676; // @[control.scala 1315:23 1512:20]
  wire [31:0] _GEN_2686 = 7'h10 == cnt_layer ? 32'h21480000 : _GEN_2677; // @[control.scala 1315:23 1513:31]
  wire [31:0] _GEN_2687 = 7'h10 == cnt_layer ? 32'h22d00000 : _GEN_2678; // @[control.scala 1315:23 1514:31]
  wire [15:0] _GEN_2688 = 7'hf == cnt_layer ? 16'h6db5 : _GEN_2679; // @[control.scala 1315:23 1495:24]
  wire [3:0] _GEN_2689 = 7'hf == cnt_layer ? 4'h8 : _GEN_2680; // @[control.scala 1315:23 1496:24]
  wire [7:0] _GEN_2690 = 7'hf == cnt_layer ? 8'h6 : _GEN_2681; // @[control.scala 1315:23 1497:19]
  wire [7:0] _GEN_2691 = 7'hf == cnt_layer ? 8'h49 : _GEN_2682; // @[control.scala 1315:23 1498:20]
  wire [31:0] _GEN_2692 = 7'hf == cnt_layer ? 32'h3e60cfdc : _GEN_2683; // @[control.scala 1315:23 1499:25]
  wire [31:0] _GEN_2693 = 7'hf == cnt_layer ? 32'h41260ba1 : _GEN_2684; // @[control.scala 1315:23 1500:25]
  wire [7:0] _GEN_2694 = 7'hf == cnt_layer ? 8'h3 : _GEN_2685; // @[control.scala 1315:23 1501:20]
  wire [31:0] _GEN_2695 = 7'hf == cnt_layer ? 32'h21438000 : _GEN_2686; // @[control.scala 1315:23 1502:31]
  wire [31:0] _GEN_2696 = 7'hf == cnt_layer ? 32'h22cff800 : _GEN_2687; // @[control.scala 1315:23 1503:31]
  wire [15:0] _GEN_2697 = 7'he == cnt_layer ? 16'h40dd : _GEN_2688; // @[control.scala 1315:23 1484:24]
  wire [3:0] _GEN_2698 = 7'he == cnt_layer ? 4'h8 : _GEN_2689; // @[control.scala 1315:23 1485:24]
  wire [7:0] _GEN_2699 = 7'he == cnt_layer ? 8'h5 : _GEN_2690; // @[control.scala 1315:23 1486:19]
  wire [7:0] _GEN_2700 = 7'he == cnt_layer ? 8'h52 : _GEN_2691; // @[control.scala 1315:23 1487:20]
  wire [31:0] _GEN_2701 = 7'he == cnt_layer ? 32'h3e01abb9 : _GEN_2692; // @[control.scala 1315:23 1488:25]
  wire [31:0] _GEN_2702 = 7'he == cnt_layer ? 32'h41a9dd98 : _GEN_2693; // @[control.scala 1315:23 1489:25]
  wire [7:0] _GEN_2703 = 7'he == cnt_layer ? 8'h6 : _GEN_2694; // @[control.scala 1315:23 1490:20]
  wire [31:0] _GEN_2704 = 7'he == cnt_layer ? 32'h213f0000 : _GEN_2695; // @[control.scala 1315:23 1491:31]
  wire [31:0] _GEN_2705 = 7'he == cnt_layer ? 32'h22cff000 : _GEN_2696; // @[control.scala 1315:23 1492:31]
  wire [15:0] _GEN_2706 = 7'hd == cnt_layer ? 16'h4198 : _GEN_2697; // @[control.scala 1315:23 1473:24]
  wire [3:0] _GEN_2707 = 7'hd == cnt_layer ? 4'h7 : _GEN_2698; // @[control.scala 1315:23 1474:24]
  wire [7:0] _GEN_2708 = 7'hd == cnt_layer ? 8'h6 : _GEN_2699; // @[control.scala 1315:23 1475:19]
  wire [7:0] _GEN_2709 = 7'hd == cnt_layer ? 8'h4a : _GEN_2700; // @[control.scala 1315:23 1476:20]
  wire [31:0] _GEN_2710 = 7'hd == cnt_layer ? 32'h3e0514bc : _GEN_2701; // @[control.scala 1315:23 1477:25]
  wire [31:0] _GEN_2711 = 7'hd == cnt_layer ? 32'h418cef57 : _GEN_2702; // @[control.scala 1315:23 1478:25]
  wire [7:0] _GEN_2712 = 7'hd == cnt_layer ? 8'h5 : _GEN_2703; // @[control.scala 1315:23 1479:20]
  wire [31:0] _GEN_2713 = 7'hd == cnt_layer ? 32'h213a8000 : _GEN_2704; // @[control.scala 1315:23 1480:31]
  wire [31:0] _GEN_2714 = 7'hd == cnt_layer ? 32'h22cfe800 : _GEN_2705; // @[control.scala 1315:23 1481:31]
  wire [15:0] _GEN_2715 = 7'hc == cnt_layer ? 16'h40b4 : _GEN_2706; // @[control.scala 1315:23 1462:24]
  wire [3:0] _GEN_2716 = 7'hc == cnt_layer ? 4'h6 : _GEN_2707; // @[control.scala 1315:23 1463:24]
  wire [7:0] _GEN_2717 = 7'hc == cnt_layer ? 8'h2 : _GEN_2708; // @[control.scala 1315:23 1464:19]
  wire [7:0] _GEN_2718 = 7'hc == cnt_layer ? 8'h4a : _GEN_2709; // @[control.scala 1315:23 1465:20]
  wire [31:0] _GEN_2719 = 7'hc == cnt_layer ? 32'h3de02dba : _GEN_2710; // @[control.scala 1315:23 1466:25]
  wire [31:0] _GEN_2720 = 7'hc == cnt_layer ? 32'h41a8091d : _GEN_2711; // @[control.scala 1315:23 1467:25]
  wire [7:0] _GEN_2721 = 7'hc == cnt_layer ? 8'h6 : _GEN_2712; // @[control.scala 1315:23 1468:20]
  wire [31:0] _GEN_2722 = 7'hc == cnt_layer ? 32'h21360000 : _GEN_2713; // @[control.scala 1315:23 1469:31]
  wire [31:0] _GEN_2723 = 7'hc == cnt_layer ? 32'h22cfe000 : _GEN_2714; // @[control.scala 1315:23 1470:31]
  wire [15:0] _GEN_2724 = 7'hb == cnt_layer ? 16'h4691 : _GEN_2715; // @[control.scala 1315:23 1451:25]
  wire [3:0] _GEN_2725 = 7'hb == cnt_layer ? 4'h7 : _GEN_2716; // @[control.scala 1315:23 1452:24]
  wire [7:0] _GEN_2726 = 7'hb == cnt_layer ? 8'h4 : _GEN_2717; // @[control.scala 1315:23 1453:19]
  wire [7:0] _GEN_2727 = 7'hb == cnt_layer ? 8'h47 : _GEN_2718; // @[control.scala 1315:23 1454:20]
  wire [31:0] _GEN_2728 = 7'hb == cnt_layer ? 32'h3e7efcb8 : _GEN_2719; // @[control.scala 1315:23 1455:25]
  wire [31:0] _GEN_2729 = 7'hb == cnt_layer ? 32'h410f6038 : _GEN_2720; // @[control.scala 1315:23 1456:25]
  wire [7:0] _GEN_2730 = 7'hb == cnt_layer ? 8'h2 : _GEN_2721; // @[control.scala 1315:23 1457:20]
  wire [31:0] _GEN_2731 = 7'hb == cnt_layer ? 32'h21318000 : _GEN_2722; // @[control.scala 1315:23 1458:31]
  wire [31:0] _GEN_2732 = 7'hb == cnt_layer ? 32'h22cfd800 : _GEN_2723; // @[control.scala 1315:23 1459:31]
  wire [15:0] _GEN_2733 = 7'ha == cnt_layer ? 16'h4f9b : _GEN_2724; // @[control.scala 1315:23 1439:25]
  wire [3:0] _GEN_2734 = 7'ha == cnt_layer ? 4'h8 : _GEN_2725; // @[control.scala 1315:23 1440:25]
  wire [7:0] _GEN_2735 = 7'ha == cnt_layer ? 8'h2 : _GEN_2726; // @[control.scala 1315:23 1441:25]
  wire [7:0] _GEN_2736 = 7'ha == cnt_layer ? 8'h5e : _GEN_2727; // @[control.scala 1315:23 1442:25]
  wire [31:0] _GEN_2737 = 7'ha == cnt_layer ? 32'h3e87cdab : _GEN_2728; // @[control.scala 1315:23 1443:25]
  wire [31:0] _GEN_2738 = 7'ha == cnt_layer ? 32'h415e7902 : _GEN_2729; // @[control.scala 1315:23 1444:25]
  wire [7:0] _GEN_2739 = 7'ha == cnt_layer ? 8'h4 : _GEN_2730; // @[control.scala 1315:23 1445:25]
  wire [31:0] _GEN_2740 = 7'ha == cnt_layer ? 32'h212d0000 : _GEN_2731; // @[control.scala 1315:23 1446:31]
  wire [31:0] _GEN_2741 = 7'ha == cnt_layer ? 32'h22cfd000 : _GEN_2732; // @[control.scala 1315:23 1447:31]
  wire [15:0] _GEN_2742 = 7'h9 == cnt_layer ? 16'h6a91 : _GEN_2733; // @[control.scala 1315:23 1426:25]
  wire [3:0] _GEN_2743 = 7'h9 == cnt_layer ? 4'h7 : _GEN_2734; // @[control.scala 1315:23 1427:25]
  wire [7:0] _GEN_2744 = 7'h9 == cnt_layer ? 8'h1 : _GEN_2735; // @[control.scala 1315:23 1428:25]
  wire [7:0] _GEN_2745 = 7'h9 == cnt_layer ? 8'h4e : _GEN_2736; // @[control.scala 1315:23 1429:25]
  wire [31:0] _GEN_2746 = 7'h9 == cnt_layer ? 32'h3ed8417b : _GEN_2737; // @[control.scala 1315:23 1430:25]
  wire [31:0] _GEN_2747 = 7'h9 == cnt_layer ? 32'h40c1d668 : _GEN_2738; // @[control.scala 1315:23 1431:25]
  wire [7:0] _GEN_2748 = 7'h9 == cnt_layer ? 8'h2 : _GEN_2739; // @[control.scala 1315:23 1432:25]
  wire [31:0] _GEN_2749 = 7'h9 == cnt_layer ? 32'h21288000 : _GEN_2740; // @[control.scala 1315:23 1433:31]
  wire [31:0] _GEN_2750 = 7'h9 == cnt_layer ? 32'h22cfc800 : _GEN_2741; // @[control.scala 1315:23 1434:31]
  wire [15:0] _GEN_2751 = 7'h8 == cnt_layer ? 16'h1 : _GEN_2742; // @[control.scala 1315:23 1415:25]
  wire [3:0] _GEN_2752 = 7'h8 == cnt_layer ? 4'h0 : _GEN_2743; // @[control.scala 1315:23 1416:25]
  wire [7:0] _GEN_2753 = 7'h8 == cnt_layer ? 8'h0 : _GEN_2744; // @[control.scala 1315:23 1417:25]
  wire [7:0] _GEN_2754 = 7'h8 == cnt_layer ? 8'h0 : _GEN_2745; // @[control.scala 1315:23 1418:25]
  wire [31:0] _GEN_2755 = 7'h8 == cnt_layer ? 32'h3f800000 : _GEN_2746; // @[control.scala 1315:23 1419:25]
  wire [31:0] _GEN_2756 = 7'h8 == cnt_layer ? 32'h3f800000 : _GEN_2747; // @[control.scala 1315:23 1420:25]
  wire [7:0] _GEN_2757 = 7'h8 == cnt_layer ? 8'h0 : _GEN_2748; // @[control.scala 1315:23 1421:25]
  wire [31:0] _GEN_2758 = 7'h8 == cnt_layer ? 32'h21240000 : _GEN_2749; // @[control.scala 1315:23 1422:31]
  wire [31:0] _GEN_2759 = 7'h8 == cnt_layer ? 32'h22cfc000 : _GEN_2750; // @[control.scala 1315:23 1423:31]
  wire [15:0] _GEN_2760 = 7'h7 == cnt_layer ? 16'h1 : _GEN_2751; // @[control.scala 1315:23 1404:25]
  wire [3:0] _GEN_2761 = 7'h7 == cnt_layer ? 4'h0 : _GEN_2752; // @[control.scala 1315:23 1405:25]
  wire [7:0] _GEN_2762 = 7'h7 == cnt_layer ? 8'h0 : _GEN_2753; // @[control.scala 1315:23 1406:25]
  wire [7:0] _GEN_2763 = 7'h7 == cnt_layer ? 8'h0 : _GEN_2754; // @[control.scala 1315:23 1407:25]
  wire [31:0] _GEN_2764 = 7'h7 == cnt_layer ? 32'h3f800000 : _GEN_2755; // @[control.scala 1315:23 1408:25]
  wire [31:0] _GEN_2765 = 7'h7 == cnt_layer ? 32'h3f800000 : _GEN_2756; // @[control.scala 1315:23 1409:25]
  wire [7:0] _GEN_2766 = 7'h7 == cnt_layer ? 8'h0 : _GEN_2757; // @[control.scala 1315:23 1410:25]
  wire [31:0] _GEN_2767 = 7'h7 == cnt_layer ? 32'h211f8000 : _GEN_2758; // @[control.scala 1315:23 1411:31]
  wire [31:0] _GEN_2768 = 7'h7 == cnt_layer ? 32'h22cfb800 : _GEN_2759; // @[control.scala 1315:23 1412:31]
  wire [15:0] _GEN_2769 = 7'h6 == cnt_layer ? 16'h1 : _GEN_2760; // @[control.scala 1315:23 1393:25]
  wire [3:0] _GEN_2770 = 7'h6 == cnt_layer ? 4'h0 : _GEN_2761; // @[control.scala 1315:23 1394:25]
  wire [7:0] _GEN_2771 = 7'h6 == cnt_layer ? 8'h0 : _GEN_2762; // @[control.scala 1315:23 1395:25]
  wire [7:0] _GEN_2772 = 7'h6 == cnt_layer ? 8'h0 : _GEN_2763; // @[control.scala 1315:23 1396:25]
  wire [31:0] _GEN_2773 = 7'h6 == cnt_layer ? 32'h3f800000 : _GEN_2764; // @[control.scala 1315:23 1397:25]
  wire [31:0] _GEN_2774 = 7'h6 == cnt_layer ? 32'h3f800000 : _GEN_2765; // @[control.scala 1315:23 1398:25]
  wire [7:0] _GEN_2775 = 7'h6 == cnt_layer ? 8'h0 : _GEN_2766; // @[control.scala 1315:23 1399:25]
  wire [31:0] _GEN_2776 = 7'h6 == cnt_layer ? 32'h211b0000 : _GEN_2767; // @[control.scala 1315:23 1400:31]
  wire [31:0] _GEN_2777 = 7'h6 == cnt_layer ? 32'h22cfb000 : _GEN_2768; // @[control.scala 1315:23 1401:31]
  wire [15:0] _GEN_2778 = 7'h5 == cnt_layer ? 16'h1 : _GEN_2769; // @[control.scala 1315:23 1382:25]
  wire [3:0] _GEN_2779 = 7'h5 == cnt_layer ? 4'h0 : _GEN_2770; // @[control.scala 1315:23 1383:25]
  wire [7:0] _GEN_2780 = 7'h5 == cnt_layer ? 8'h0 : _GEN_2771; // @[control.scala 1315:23 1384:25]
  wire [7:0] _GEN_2781 = 7'h5 == cnt_layer ? 8'h0 : _GEN_2772; // @[control.scala 1315:23 1385:25]
  wire [31:0] _GEN_2782 = 7'h5 == cnt_layer ? 32'h3f800000 : _GEN_2773; // @[control.scala 1315:23 1386:25]
  wire [31:0] _GEN_2783 = 7'h5 == cnt_layer ? 32'h3f800000 : _GEN_2774; // @[control.scala 1315:23 1387:25]
  wire [7:0] _GEN_2784 = 7'h5 == cnt_layer ? 8'h0 : _GEN_2775; // @[control.scala 1315:23 1388:25]
  wire [31:0] _GEN_2785 = 7'h5 == cnt_layer ? 32'h21168000 : _GEN_2776; // @[control.scala 1315:23 1389:31]
  wire [31:0] _GEN_2786 = 7'h5 == cnt_layer ? 32'h22cfa800 : _GEN_2777; // @[control.scala 1315:23 1390:31]
  wire [15:0] _GEN_2787 = 7'h4 == cnt_layer ? 16'h78fa : _GEN_2778; // @[control.scala 1315:23 1371:25]
  wire [3:0] _GEN_2788 = 7'h4 == cnt_layer ? 4'h8 : _GEN_2779; // @[control.scala 1315:23 1372:25]
  wire [7:0] _GEN_2789 = 7'h4 == cnt_layer ? 8'h1 : _GEN_2780; // @[control.scala 1315:23 1373:25]
  wire [7:0] _GEN_2790 = 7'h4 == cnt_layer ? 8'h46 : _GEN_2781; // @[control.scala 1315:23 1374:25]
  wire [31:0] _GEN_2791 = 7'h4 == cnt_layer ? 32'h3f37d0c3 : _GEN_2782; // @[control.scala 1315:23 1375:25]
  wire [31:0] _GEN_2792 = 7'h4 == cnt_layer ? 32'h4046a036 : _GEN_2783; // @[control.scala 1315:23 1376:25]
  wire [7:0] _GEN_2793 = 7'h4 == cnt_layer ? 8'h1 : _GEN_2784; // @[control.scala 1315:23 1377:25]
  wire [31:0] _GEN_2794 = 7'h4 == cnt_layer ? 32'h21120000 : _GEN_2785; // @[control.scala 1315:23 1378:31]
  wire [31:0] _GEN_2795 = 7'h4 == cnt_layer ? 32'h22cfa000 : _GEN_2786; // @[control.scala 1315:23 1379:31]
  wire [15:0] _GEN_2796 = 7'h3 == cnt_layer ? 16'h601d : _GEN_2787; // @[control.scala 1315:23 1360:25]
  wire [3:0] _GEN_2797 = 7'h3 == cnt_layer ? 4'h6 : _GEN_2788; // @[control.scala 1315:23 1361:25]
  wire [7:0] _GEN_2798 = 7'h3 == cnt_layer ? 8'h1 : _GEN_2789; // @[control.scala 1315:23 1362:25]
  wire [7:0] _GEN_2799 = 7'h3 == cnt_layer ? 8'h42 : _GEN_2790; // @[control.scala 1315:23 1363:25]
  wire [31:0] _GEN_2800 = 7'h3 == cnt_layer ? 32'h3f45347f : _GEN_2791; // @[control.scala 1315:23 1364:25]
  wire [31:0] _GEN_2801 = 7'h3 == cnt_layer ? 32'h402c147b : _GEN_2792; // @[control.scala 1315:23 1365:25]
  wire [7:0] _GEN_2802 = 7'h3 == cnt_layer ? 8'h1 : _GEN_2793; // @[control.scala 1315:23 1366:25]
  wire [31:0] _GEN_2803 = 7'h3 == cnt_layer ? 32'h210d8000 : _GEN_2794; // @[control.scala 1315:23 1367:31]
  wire [31:0] _GEN_2804 = 7'h3 == cnt_layer ? 32'h22cf9800 : _GEN_2795; // @[control.scala 1315:23 1368:31]
  wire [25:0] _GEN_2860 = reset ? 26'h0 : _GEN_1899; // @[control.scala 180:{34,34}]
  wire [34:0] _GEN_2861 = reset ? 35'h0 : _ifm_addr_t_T_2; // @[control.scala 380:{29,29} 413:16]
  wire [34:0] _GEN_2862 = reset ? 35'h0 : _ofm_addr_t_T_2; // @[control.scala 415:{29,29} 417:16]
  wire [9:0] _GEN_2863 = reset ? 10'h0 : _GEN_1890; // @[control.scala 425:{46,46}]
  assign io_conv_finish = conv_finish; // @[control.scala 72:19]
  assign io_reg0 = reg_t_0; // @[control.scala 166:12]
  assign io_reg1 = reg_t_1; // @[control.scala 167:12]
  assign io_reg2 = reg_t_2; // @[control.scala 168:12]
  assign io_reg3 = reg_t_3; // @[control.scala 169:12]
  assign io_reg4 = reg_t_4; // @[control.scala 170:12]
  assign io_reg5 = reg_t_5; // @[control.scala 171:12]
  assign io_reg6 = reg_t_6; // @[control.scala 172:12]
  assign io_reg7 = reg_t_7; // @[control.scala 173:12]
  assign io_reg8 = reg_t_8; // @[control.scala 174:12]
  assign io_reg9 = reg_t_9; // @[control.scala 175:12]
  assign io_reg10 = reg_t_10; // @[control.scala 176:13]
  assign io_yolo_finish = ~io_yolo_finish_REG & yolo_finish; // @[utils.scala 10:27]
  assign io_resize_load = resize_load_t; // @[control.scala 421:20]
  always @(posedge clock) begin
    if (reset) begin // @[control.scala 40:28]
      yolo_finish <= 1'h0; // @[control.scala 40:28]
    end else if (6'h0 == state) begin // @[control.scala 438:19]
      yolo_finish <= 1'h0; // @[control.scala 444:25]
    end else if (!(6'h1 == state)) begin // @[control.scala 438:19]
      if (!(6'h2 == state)) begin // @[control.scala 438:19]
        yolo_finish <= _GEN_1768;
      end
    end
    if (reset) begin // @[utils.scala 10:17]
      io_yolo_finish_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      io_yolo_finish_REG <= yolo_finish; // @[utils.scala 10:17]
    end
    if (reset) begin // @[utils.scala 10:17]
      ap_done_up_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      ap_done_up_REG <= io_ap_done; // @[utils.scala 10:17]
    end
    if (reset) begin // @[control.scala 46:26]
      c2f_cnt <= 4'h0; // @[control.scala 46:26]
    end else if (current_layer != current_layer_next & current_layer_is_c2f_next) begin // @[control.scala 85:19]
      if (_c2f_shortcut_T_6) begin // @[control.scala 85:91]
        c2f_cnt <= 4'h0;
      end else begin
        c2f_cnt <= _c2f_cnt_T_4;
      end
    end
    if (reset) begin // @[control.scala 52:32]
      current_layer <= 5'h0; // @[control.scala 52:32]
    end else if (layer_finish) begin // @[control.scala 109:25]
      if (cur_layer_sel_21) begin // @[control.scala 109:43]
        current_layer <= 5'h0;
      end else begin
        current_layer <= _current_layer_T_2;
      end
    end
    if (reset) begin // @[control.scala 71:30]
      conv_finish <= 1'h0; // @[control.scala 71:30]
    end else if (6'h0 == state) begin // @[control.scala 438:19]
      conv_finish <= 1'h0; // @[control.scala 443:25]
    end else if (!(6'h1 == state)) begin // @[control.scala 438:19]
      if (!(6'h2 == state)) begin // @[control.scala 438:19]
        conv_finish <= _GEN_1769;
      end
    end
    current_layer_next <= current_layer; // @[control.scala 81:37]
    current_layer_is_c2f_next <= current_model_code == 3'h1; // @[control.scala 76:51]
    if (reset) begin // @[control.scala 90:34]
      conv_cnt_in_c2f <= 5'h0; // @[control.scala 90:34]
    end else if (current_layer_is_c2f & conv_finish) begin // @[control.scala 91:27]
      if (conv_cnt_in_c2f == _conv_cnt_in_c2f_T_2) begin // @[control.scala 91:67]
        conv_cnt_in_c2f <= 5'h0;
      end else begin
        conv_cnt_in_c2f <= _conv_cnt_in_c2f_T_5;
      end
    end
    if (reset) begin // @[control.scala 93:30]
      cnt_in_sppf <= 3'h0; // @[control.scala 93:30]
    end else if (current_layer_is_sppf & conv_finish) begin // @[control.scala 94:23]
      if (cnt_in_sppf == 3'h1) begin // @[control.scala 94:64]
        cnt_in_sppf <= 3'h0;
      end else begin
        cnt_in_sppf <= _cnt_in_sppf_T_3;
      end
    end
    if (reset) begin // @[control.scala 96:36]
      cnt_in_detect_box <= 3'h0; // @[control.scala 96:36]
    end else if (current_layer_is_detect_box & conv_finish) begin // @[control.scala 97:29]
      if (cnt_in_detect_box == 3'h2) begin // @[control.scala 97:76]
        cnt_in_detect_box <= 3'h0;
      end else begin
        cnt_in_detect_box <= _cnt_in_detect_box_T_3;
      end
    end
    if (reset) begin // @[control.scala 99:36]
      cnt_in_detect_cls <= 3'h0; // @[control.scala 99:36]
    end else if (current_layer_is_detect_cls & conv_finish) begin // @[control.scala 100:29]
      if (cnt_in_detect_cls == 3'h2) begin // @[control.scala 100:76]
        cnt_in_detect_cls <= 3'h0;
      end else begin
        cnt_in_detect_cls <= _cnt_in_detect_cls_T_3;
      end
    end
    if (reset) begin // @[control.scala 112:28]
      conv_scale <= 16'h0; // @[control.scala 112:28]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      conv_scale <= 16'h4741; // @[control.scala 1320:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      conv_scale <= 16'h44b7; // @[control.scala 1333:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      conv_scale <= 16'h5116; // @[control.scala 1349:25]
    end else begin
      conv_scale <= _GEN_2796;
    end
    if (reset) begin // @[control.scala 113:29]
      conv_shift <= 4'h0; // @[control.scala 113:29]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      conv_shift <= 4'h9; // @[control.scala 1321:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      conv_shift <= 4'h7; // @[control.scala 1334:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      conv_shift <= 4'h6; // @[control.scala 1350:25]
    end else begin
      conv_shift <= _GEN_2797;
    end
    if (reset) begin // @[control.scala 114:24]
      zp_in <= 8'h0; // @[control.scala 114:24]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      zp_in <= 8'h0; // @[control.scala 1322:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      zp_in <= 8'h1; // @[control.scala 1335:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      zp_in <= 8'h0; // @[control.scala 1351:25]
    end else begin
      zp_in <= _GEN_2798;
    end
    if (reset) begin // @[control.scala 115:25]
      zp_out <= 8'h0; // @[control.scala 115:25]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      zp_out <= 8'h41; // @[control.scala 1323:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      zp_out <= 8'h3d; // @[control.scala 1336:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      zp_out <= 8'h5b; // @[control.scala 1352:25]
    end else begin
      zp_out <= _GEN_2799;
    end
    if (reset) begin // @[control.scala 116:25]
      zp_act <= 8'h0; // @[control.scala 116:25]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      zp_act <= 8'h1; // @[control.scala 1326:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      zp_act <= 8'h0; // @[control.scala 1339:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      zp_act <= 8'h1; // @[control.scala 1355:25]
    end else begin
      zp_act <= _GEN_2802;
    end
    if (reset) begin // @[control.scala 117:30]
      scale_B_act <= 32'h0; // @[control.scala 117:30]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      scale_B_act <= 32'h3f7e6443; // @[control.scala 1324:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      scale_B_act <= 32'h402c4204; // @[control.scala 1337:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      scale_B_act <= 32'h3faedda2; // @[control.scala 1353:25]
    end else begin
      scale_B_act <= _GEN_2800;
    end
    if (reset) begin // @[control.scala 118:30]
      scale_A_act <= 32'h0; // @[control.scala 118:30]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      scale_A_act <= 32'h4003061c; // @[control.scala 1325:25]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      scale_A_act <= 32'h3f3668c2; // @[control.scala 1338:25]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      scale_A_act <= 32'h4025ea3b; // @[control.scala 1354:25]
    end else begin
      scale_A_act <= _GEN_2801;
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_0 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        reg_t_0 <= 32'h209; // @[control.scala 475:22]
      end else if (6'h2 == state) begin // @[control.scala 438:19]
        reg_t_0 <= _GEN_7;
      end else begin
        reg_t_0 <= _GEN_1728;
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_1 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_1 <= _GEN_1730;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_2 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_2 <= _GEN_1731;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_3 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_3 <= _GEN_1742;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_4 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        reg_t_4 <= bia_ddr_base_addr; // @[control.scala 473:22]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        reg_t_4 <= _GEN_1726;
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_5 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        reg_t_5 <= {{13'd0}, _reg_t_5_T}; // @[control.scala 474:22]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        reg_t_5 <= _GEN_1727;
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_6 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_6 <= _GEN_1763;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_7 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_7 <= _GEN_1764;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_8 <= 32'h0; // @[control.scala 160:37]
    end else begin
      reg_t_8 <= _reg_t_8_T_1; // @[control.scala 306:14]
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_9 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_9 <= _GEN_1732;
        end
      end
    end
    if (reset) begin // @[control.scala 160:37]
      reg_t_10 <= 32'h0; // @[control.scala 160:37]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_t_10 <= _GEN_1733;
        end
      end
    end
    if (reset) begin // @[control.scala 161:29]
      reg_static <= 32'h0; // @[control.scala 161:29]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_static <= _GEN_1739;
        end
      end
    end
    if (reset) begin // @[control.scala 162:27]
      reg_task <= 32'h0; // @[control.scala 162:27]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          reg_task <= _GEN_1741;
        end
      end
    end
    if (reset) begin // @[control.scala 163:24]
      cnt_t <= 5'h0; // @[control.scala 163:24]
    end else if (6'h0 == state) begin // @[control.scala 438:19]
      cnt_t <= _GEN_2;
    end else if (6'h1 == state) begin // @[control.scala 438:19]
      cnt_t <= 5'h0; // @[control.scala 476:19]
    end else if (6'h2 == state) begin // @[control.scala 438:19]
      cnt_t <= _GEN_2;
    end else begin
      cnt_t <= _GEN_1729;
    end
    if (reset) begin // @[control.scala 178:32]
      wgt_addr_send <= 32'h0; // @[control.scala 178:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        wgt_addr_send <= wgt_ddr_base_addr; // @[control.scala 462:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        wgt_addr_send <= _GEN_1751;
      end
    end
    if (reset) begin // @[control.scala 179:32]
      wgt_addr_read <= 16'h0; // @[control.scala 179:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        wgt_addr_read <= 16'h0; // @[control.scala 463:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        wgt_addr_read <= _GEN_1752;
      end
    end
    wgt_addr_read_t <= _GEN_2860[15:0]; // @[control.scala 180:{34,34}]
    if (reset) begin // @[control.scala 181:32]
      bia_addr_read <= 16'h0; // @[control.scala 181:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        bia_addr_read <= 16'h0; // @[control.scala 464:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        bia_addr_read <= _GEN_1761;
      end
    end
    if (reset) begin // @[control.scala 182:31]
      last_buf_sel <= 1'h0; // @[control.scala 182:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        last_buf_sel <= 1'h0; // @[control.scala 465:26]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        last_buf_sel <= _GEN_1740;
      end
    end
    if (reset) begin // @[control.scala 192:31]
      iter_ifm_pre <= 13'h0; // @[control.scala 192:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_ifm_pre <= 13'h0; // @[control.scala 466:26]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_ifm_pre <= _GEN_1756;
      end
    end
    if (reset) begin // @[control.scala 194:31]
      iter_ofm_pre <= 13'h0; // @[control.scala 194:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_ofm_pre <= 13'h0; // @[control.scala 467:26]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_ofm_pre <= _GEN_1758;
      end
    end
    if (reset) begin // @[control.scala 195:31]
      iter_div_pre <= 13'h0; // @[control.scala 195:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_div_pre <= 13'h0; // @[control.scala 468:26]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_div_pre <= _GEN_1757;
      end
    end
    if (reset) begin // @[control.scala 196:32]
      iter_ifm_post <= 13'h0; // @[control.scala 196:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_ifm_post <= 13'h0; // @[control.scala 469:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_ifm_post <= _GEN_1753;
      end
    end
    if (reset) begin // @[control.scala 197:32]
      iter_ofm_post <= 13'h0; // @[control.scala 197:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_ofm_post <= 13'h0; // @[control.scala 470:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_ofm_post <= _GEN_1755;
      end
    end
    if (reset) begin // @[control.scala 198:32]
      iter_div_post <= 13'h0; // @[control.scala 198:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        iter_div_post <= 13'h0; // @[control.scala 471:27]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        iter_div_post <= _GEN_1754;
      end
    end
    if (reset) begin // @[control.scala 274:27]
      weight_sel <= 3'h0; // @[control.scala 274:27]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          weight_sel <= _GEN_1760;
        end
      end
    end
    if (reset) begin // @[control.scala 290:27]
      pool_cnt <= 2'h0; // @[control.scala 290:27]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        pool_cnt <= 2'h0; // @[control.scala 461:21]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        pool_cnt <= _GEN_1765;
      end
    end
    if (reset) begin // @[control.scala 295:38]
      bottleneck_transfer <= 1'h0; // @[control.scala 295:38]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        bottleneck_transfer <= 1'h0; // @[control.scala 459:33]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        bottleneck_transfer <= _GEN_1743;
      end
    end
    if (reset) begin // @[control.scala 296:35]
      bottleneck_ready <= 1'h0; // @[control.scala 296:35]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        bottleneck_ready <= 1'h0; // @[control.scala 460:30]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        bottleneck_ready <= _GEN_1744;
      end
    end
    if (reset) begin // @[control.scala 299:33]
      cnt_detect_cls <= 2'h0; // @[control.scala 299:33]
    end else if (_c2f_cnt_T & current_layer_is_detect_cls_next) begin // @[control.scala 301:26]
      if (cnt_detect_cls == 2'h2) begin // @[control.scala 301:105]
        cnt_detect_cls <= 2'h0;
      end else begin
        cnt_detect_cls <= _cnt_detect_cls_T_4;
      end
    end
    current_layer_is_detect_cls_next <= current_model_code == 3'h4; // @[control.scala 79:58]
    if (reset) begin // @[control.scala 316:41]
      iter_div_prexfm_div_col <= 32'h0; // @[control.scala 316:41]
    end else begin
      iter_div_prexfm_div_col <= {{4'd0}, _iter_div_prexfm_div_col_T}; // @[control.scala 332:29]
    end
    if (reset) begin // @[control.scala 319:41]
      fm_row_fm_res_t1xfm_col <= 32'h0; // @[control.scala 319:41]
    end else begin
      fm_row_fm_res_t1xfm_col <= {{12'd0}, _fm_row_fm_res_t1xfm_col_T_2}; // @[control.scala 334:28]
    end
    if (reset) begin // @[control.scala 320:38]
      fm_row_fm_resxfm_col <= 32'h0; // @[control.scala 320:38]
    end else begin
      fm_row_fm_resxfm_col <= {{12'd0}, _fm_row_fm_resxfm_col_T_2}; // @[control.scala 335:25]
    end
    if (reset) begin // @[control.scala 352:44]
      iter_div_postxfm_col_output <= 32'h0; // @[control.scala 352:44]
    end else begin
      iter_div_postxfm_col_output <= {{3'd0}, _iter_div_postxfm_col_output_T_1}; // @[control.scala 354:32]
    end
    if (reset) begin // @[control.scala 353:48]
      fm_row_res_outputxfm_col_output <= 32'h0; // @[control.scala 353:48]
    end else begin
      fm_row_res_outputxfm_col_output <= {{12'd0}, _fm_row_res_outputxfm_col_output_T_2}; // @[control.scala 355:36]
    end
    if (reset) begin // @[control.scala 357:39]
      ifm_send_task_enable <= 1'h0; // @[control.scala 357:39]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ifm_send_task_enable <= _GEN_1734;
        end
      end
    end
    if (reset) begin // @[control.scala 358:39]
      ofm_recv_task_enable <= 1'h0; // @[control.scala 358:39]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ofm_recv_task_enable <= _GEN_1745;
        end
      end
    end
    if (reset) begin // @[control.scala 359:39]
      wgt_send_task_enable <= 1'h0; // @[control.scala 359:39]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          wgt_send_task_enable <= _GEN_1750;
        end
      end
    end
    if (reset) begin // @[control.scala 362:34]
      ifm_addr_fmbase <= 32'h0; // @[control.scala 362:34]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ifm_addr_fmbase <= _GEN_1735;
        end
      end
    end
    if (reset) begin // @[control.scala 363:34]
      ifm_addr_offset <= 32'h0; // @[control.scala 363:34]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ifm_addr_offset <= _GEN_1736;
        end
      end
    end
    if (reset) begin // @[control.scala 364:31]
      ifm_send_len <= 32'h0; // @[control.scala 364:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ifm_send_len <= _GEN_1737;
        end
      end
    end
    if (reset) begin // @[control.scala 365:34]
      ofm_addr_fmbase <= 32'h0; // @[control.scala 365:34]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ofm_addr_fmbase <= _GEN_1747;
        end
      end
    end
    if (reset) begin // @[control.scala 366:34]
      ofm_addr_offset <= 32'h0; // @[control.scala 366:34]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ofm_addr_offset <= _GEN_1748;
        end
      end
    end
    if (reset) begin // @[control.scala 367:31]
      ofm_recv_len <= 32'h0; // @[control.scala 367:31]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ofm_recv_len <= _GEN_1749;
        end
      end
    end
    if (reset) begin // @[control.scala 369:36]
      wgt_ddr_base_addr <= 32'h0; // @[control.scala 369:36]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      wgt_ddr_base_addr <= 32'h21000000; // @[control.scala 1327:31]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      wgt_ddr_base_addr <= 32'h21048000; // @[control.scala 1340:31]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      wgt_ddr_base_addr <= 32'h21090000; // @[control.scala 1356:31]
    end else begin
      wgt_ddr_base_addr <= _GEN_2803;
    end
    if (reset) begin // @[control.scala 370:36]
      bia_ddr_base_addr <= 32'h0; // @[control.scala 370:36]
    end else if (7'h0 == cnt_layer) begin // @[control.scala 1315:23]
      bia_ddr_base_addr <= 32'h22cf8000; // @[control.scala 1328:31]
    end else if (7'h1 == cnt_layer) begin // @[control.scala 1315:23]
      bia_ddr_base_addr <= 32'h22cf8800; // @[control.scala 1341:31]
    end else if (7'h2 == cnt_layer) begin // @[control.scala 1315:23]
      bia_ddr_base_addr <= 32'h22cf9000; // @[control.scala 1357:31]
    end else begin
      bia_ddr_base_addr <= _GEN_2804;
    end
    if (reset) begin // @[control.scala 379:24]
      ifm_sel <= 1'h0; // @[control.scala 379:24]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          ifm_sel <= _GEN_1766;
        end
      end
    end
    ifm_addr_t <= _GEN_2861[31:0]; // @[control.scala 380:{29,29} 413:16]
    if (reset) begin // @[control.scala 381:32]
      ifm_addr_send <= 32'h0; // @[control.scala 381:32]
    end else begin
      ifm_addr_send <= _ifm_addr_send_T_2; // @[control.scala 414:19]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ifm_ddr_base_addr_regnext1 <= 32'h0; // @[Reg.scala 35:20]
    end else if (conv_finish) begin // @[Reg.scala 36:18]
      if (current_layer_is_conv | _upsample_en_T_1 | pool_en | current_layer_is_detect_cls & cnt_in_detect_cls == 3'h0
         | current_layer_is_detect_box & cnt_in_detect_box == 3'h0) begin // @[control.scala 408:29]
        if (5'h15 == current_layer) begin // @[Mux.scala 81:58]
          ifm_ddr_base_addr_regnext1 <= 32'h20e4e800;
        end else begin
          ifm_ddr_base_addr_regnext1 <= _ifm_ddr_base_addr_t_T_41;
        end
      end else if (current_layer_is_c2f) begin // @[control.scala 405:34]
        ifm_ddr_base_addr_regnext1 <= ifm_ddr_base_addr_temp_c2f;
      end else begin
        ifm_ddr_base_addr_regnext1 <= _ifm_ddr_base_addr_temp_T;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      ifm_ddr_base_addr_regnext2 <= 32'h0; // @[Reg.scala 35:20]
    end else if (conv_finish) begin // @[Reg.scala 36:18]
      ifm_ddr_base_addr_regnext2 <= ifm_ddr_base_addr_regnext1; // @[Reg.scala 36:22]
    end
    ofm_addr_t <= _GEN_2862[31:0]; // @[control.scala 415:{29,29} 417:16]
    if (reset) begin // @[control.scala 416:32]
      ofm_addr_recv <= 32'h0; // @[control.scala 416:32]
    end else begin
      ofm_addr_recv <= _ofm_addr_recv_T_1; // @[control.scala 418:19]
    end
    if (reset) begin // @[control.scala 420:32]
      resize_load_t <= 1'h0; // @[control.scala 420:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (!(6'h1 == state)) begin // @[control.scala 438:19]
        if (!(6'h2 == state)) begin // @[control.scala 438:19]
          resize_load_t <= _GEN_1767;
        end
      end
    end
    if (reset) begin // @[control.scala 422:38]
      first_ofm_recv_stop <= 1'h0; // @[control.scala 422:38]
    end else if (6'h0 == state) begin // @[control.scala 438:19]
      first_ofm_recv_stop <= cur_layer_sel_0;
    end else if (!(6'h1 == state)) begin // @[control.scala 438:19]
      if (!(6'h2 == state)) begin // @[control.scala 438:19]
        first_ofm_recv_stop <= _GEN_1746;
      end
    end
    if (reset) begin // @[control.scala 424:32]
      wgt_ddr_read_en <= 1'h0; // @[control.scala 424:32]
    end else if (!(6'h0 == state)) begin // @[control.scala 438:19]
      if (6'h1 == state) begin // @[control.scala 438:19]
        wgt_ddr_read_en <= 1'h0; // @[control.scala 472:28]
      end else if (!(6'h2 == state)) begin // @[control.scala 438:19]
        wgt_ddr_read_en <= _GEN_1762;
      end
    end
    the_number_of_row_transferred <= _GEN_2863[7:0]; // @[control.scala 425:{46,46}]
    if (reset) begin // @[control.scala 436:24]
      state <= 6'h0; // @[control.scala 436:24]
    end else if (6'h0 == state) begin // @[control.scala 438:19]
      if (cnt_t_is_5) begin // @[control.scala 445:30]
        state <= 6'h1; // @[control.scala 447:23]
      end
    end else if (6'h1 == state) begin // @[control.scala 438:19]
      state <= 6'h2; // @[control.scala 477:19]
    end else if (6'h2 == state) begin // @[control.scala 438:19]
      state <= _GEN_6;
    end else begin
      state <= _GEN_1725;
    end
    if (reset) begin // @[control.scala 1305:25]
      conv_cnt <= 1'h0; // @[control.scala 1305:25]
    end else if (layer_finish) begin // @[control.scala 1308:18]
      conv_cnt <= 1'h0;
    end else if (conv_finish) begin // @[control.scala 1308:39]
      conv_cnt <= conv_cnt + 1'h1;
    end
    if (reset) begin // @[control.scala 1309:21]
      base <= 7'h0; // @[control.scala 1309:21]
    end else if (layer_finish) begin // @[control.scala 1313:14]
      if (cur_layer_sel_21) begin // @[control.scala 1313:31]
        base <= 7'h0;
      end else begin
        base <= _base_T_2;
      end
    end
    if (reset) begin // @[control.scala 1312:28]
      cnt_layer <= 7'h0; // @[control.scala 1312:28]
    end else begin
      cnt_layer <= _cnt_layer_T_1; // @[control.scala 1314:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  yolo_finish = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_yolo_finish_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ap_done_up_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  c2f_cnt = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  current_layer = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  conv_finish = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  current_layer_next = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  current_layer_is_c2f_next = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  conv_cnt_in_c2f = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  cnt_in_sppf = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  cnt_in_detect_box = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  cnt_in_detect_cls = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  conv_scale = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  conv_shift = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  zp_in = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  zp_out = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  zp_act = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  scale_B_act = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  scale_A_act = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  reg_t_0 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  reg_t_1 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg_t_2 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg_t_3 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg_t_4 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  reg_t_5 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  reg_t_6 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  reg_t_7 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  reg_t_8 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  reg_t_9 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  reg_t_10 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  reg_static = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  reg_task = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  cnt_t = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  wgt_addr_send = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  wgt_addr_read = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  wgt_addr_read_t = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  bia_addr_read = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  last_buf_sel = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  iter_ifm_pre = _RAND_38[12:0];
  _RAND_39 = {1{`RANDOM}};
  iter_ofm_pre = _RAND_39[12:0];
  _RAND_40 = {1{`RANDOM}};
  iter_div_pre = _RAND_40[12:0];
  _RAND_41 = {1{`RANDOM}};
  iter_ifm_post = _RAND_41[12:0];
  _RAND_42 = {1{`RANDOM}};
  iter_ofm_post = _RAND_42[12:0];
  _RAND_43 = {1{`RANDOM}};
  iter_div_post = _RAND_43[12:0];
  _RAND_44 = {1{`RANDOM}};
  weight_sel = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  pool_cnt = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  bottleneck_transfer = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  bottleneck_ready = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  cnt_detect_cls = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  current_layer_is_detect_cls_next = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  iter_div_prexfm_div_col = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  fm_row_fm_res_t1xfm_col = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  fm_row_fm_resxfm_col = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  iter_div_postxfm_col_output = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  fm_row_res_outputxfm_col_output = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  ifm_send_task_enable = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ofm_recv_task_enable = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  wgt_send_task_enable = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  ifm_addr_fmbase = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  ifm_addr_offset = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  ifm_send_len = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  ofm_addr_fmbase = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  ofm_addr_offset = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  ofm_recv_len = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  wgt_ddr_base_addr = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  bia_ddr_base_addr = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  ifm_sel = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  ifm_addr_t = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  ifm_addr_send = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  ifm_ddr_base_addr_regnext1 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  ifm_ddr_base_addr_regnext2 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  ofm_addr_t = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  ofm_addr_recv = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  resize_load_t = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  first_ofm_recv_stop = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  wgt_ddr_read_en = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  the_number_of_row_transferred = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  state = _RAND_77[5:0];
  _RAND_78 = {1{`RANDOM}};
  conv_cnt = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  base = _RAND_79[6:0];
  _RAND_80 = {1{`RANDOM}};
  cnt_layer = _RAND_80[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module control_signal(
  input         clock,
  input         reset,
  input         io_shutdown,
  input         io_skip_act,
  input  [9:0]  io_conv_col,
  input  [9:0]  io_conv_row,
  input         io_s_mod,
  input         io_kernal,
  output [10:0] io_ifmbuf_bram_addr_read_s1,
  output        io_ifmbuf_addr_read_sel_s1,
  output [9:0]  io_ifmbuf_bram_addr_read_s2_singal,
  output [9:0]  io_ifmbuf_bram_addr_read_s2_double,
  output [11:0] io_acc_read_addr,
  output [11:0] io_acc_write_addr,
  output        io_acc_read_en,
  output        io_acc_write_en,
  output        io_acc_curr_data_zero,
  output [11:0] io_ofm_addr,
  output        io_ofm_valid,
  output        io_ofm_done,
  input         io_pad_top,
  input         io_pad_bottom,
  input         io_pad_left_and_right,
  input         io_pad_size,
  output        io_zero_pad_valid_s1,
  output [4:0]  io_zero_pad_valid_s2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] stride = io_s_mod ? 2'h2 : 2'h1; // @[control.scala 2750:16]
  wire [1:0] _conv_col_include_pad_T = {io_pad_size, 1'h0}; // @[control.scala 2754:82]
  wire [1:0] _conv_col_include_pad_T_1 = io_pad_left_and_right ? _conv_col_include_pad_T : 2'h0; // @[control.scala 2754:46]
  wire [9:0] _GEN_131 = {{8'd0}, _conv_col_include_pad_T_1}; // @[control.scala 2754:41]
  wire [9:0] conv_col_include_pad = io_conv_col + _GEN_131; // @[control.scala 2754:41]
  wire  _conv_row_include_pad_T_1 = io_pad_bottom & io_pad_top; // @[control.scala 2755:94]
  wire [1:0] _conv_row_include_pad_T_3 = io_pad_bottom & io_pad_top ? _conv_col_include_pad_T : {{1'd0}, io_pad_size}; // @[control.scala 2755:79]
  wire [1:0] _conv_row_include_pad_T_4 = io_pad_bottom | io_pad_top ? _conv_row_include_pad_T_3 : 2'h0; // @[control.scala 2755:46]
  wire [9:0] _GEN_132 = {{8'd0}, _conv_row_include_pad_T_4}; // @[control.scala 2755:41]
  wire [9:0] conv_row_include_pad = io_conv_row + _GEN_132; // @[control.scala 2755:41]
  wire [9:0] _GEN_133 = {{8'd0}, stride}; // @[control.scala 2762:51]
  wire [9:0] conv_col_minus_stride = conv_col_include_pad - _GEN_133; // @[control.scala 2762:51]
  reg [9:0] col_cnt; // @[control.scala 2766:26]
  reg [9:0] row_cnt; // @[control.scala 2767:26]
  wire  _col_cnt_T = col_cnt == conv_col_minus_stride; // @[control.scala 2769:43]
  wire [9:0] _col_cnt_T_3 = col_cnt + _GEN_133; // @[control.scala 2769:84]
  wire [9:0] _row_cnt_T_2 = row_cnt + _GEN_133; // @[control.scala 2770:83]
  wire [9:0] _GEN_136 = {{9'd0}, io_pad_size}; // @[control.scala 2780:67]
  wire [9:0] _zero_pad_left_and_right_T_2 = io_conv_col + _GEN_136; // @[control.scala 2780:110]
  wire  zero_pad_left_and_right = io_pad_left_and_right & (col_cnt < _GEN_136 | col_cnt >= _zero_pad_left_and_right_T_2)
    ; // @[control.scala 2780:55]
  wire  zero_pad_top = io_pad_top & row_cnt < _GEN_136; // @[control.scala 2781:33]
  wire  _zero_pad_only_bottom_T_1 = io_pad_bottom & ~io_pad_top; // @[control.scala 2782:44]
  wire  zero_pad_only_bottom = io_pad_bottom & ~io_pad_top & row_cnt >= io_conv_row; // @[control.scala 2782:60]
  wire [9:0] _zero_pad_bottom_include_top_T_2 = io_conv_row + _GEN_136; // @[control.scala 2783:91]
  wire  zero_pad_bottom_include_top = _conv_row_include_pad_T_1 & row_cnt >= _zero_pad_bottom_include_top_T_2; // @[control.scala 2783:64]
  wire  zero_pad = zero_pad_left_and_right | zero_pad_top | zero_pad_bottom_include_top | zero_pad_only_bottom; // @[control.scala 2784:88]
  reg  io_zero_pad_valid_s1_REG; // @[control.scala 2785:36]
  wire  zero_s2_pad_left = io_pad_left_and_right & col_cnt == 10'h0; // @[control.scala 2792:47]
  wire  zero_s2_pad_right = io_pad_left_and_right & col_cnt == io_conv_col; // @[control.scala 2793:48]
  wire  zero_s2_pad_top = io_pad_top & row_cnt == 10'h0; // @[control.scala 2794:35]
  wire [9:0] _zero_s2_pad_only_bottom_T_3 = io_conv_row - 10'h1; // @[control.scala 2795:86]
  wire  zero_s2_pad_only_bottom = _zero_pad_only_bottom_T_1 & row_cnt == _zero_s2_pad_only_bottom_T_3; // @[control.scala 2795:60]
  wire  zero_s2_pad_bottom_include_top = _conv_row_include_pad_T_1 & row_cnt == io_conv_row; // @[control.scala 2796:67]
  wire [1:0] io_zero_pad_valid_s2_lo = {zero_s2_pad_only_bottom,zero_s2_pad_bottom_include_top}; // @[Cat.scala 33:92]
  wire [2:0] io_zero_pad_valid_s2_hi = {zero_s2_pad_left,zero_s2_pad_right,zero_s2_pad_top}; // @[Cat.scala 33:92]
  reg [4:0] io_zero_pad_valid_s2_REG; // @[control.scala 2798:35]
  reg  row_is_singal_or_double; // @[control.scala 2800:42]
  wire  _row_is_singal_or_double_T_1 = ~row_is_singal_or_double; // @[control.scala 2803:97]
  wire  _row_is_singal_T = ~zero_pad; // @[control.scala 2804:24]
  wire  _row_is_singal_T_3 = ~io_s_mod; // @[control.scala 2804:69]
  wire  _row_is_singal_T_7 = ~_col_cnt_T; // @[control.scala 2804:135]
  wire  row_is_singal = ~zero_pad & _row_is_singal_or_double_T_1 & ~io_s_mod | io_s_mod & ~
    zero_s2_pad_bottom_include_top & ~_col_cnt_T; // @[control.scala 2804:81]
  wire  row_is_double = _row_is_singal_T & row_is_singal_or_double & _row_is_singal_T_3 | io_s_mod & ~zero_s2_pad_top &
    _row_is_singal_T_7; // @[control.scala 2805:78]
  reg [10:0] bram_read_addr_singal; // @[control.scala 2807:40]
  reg [10:0] bram_read_addr_double; // @[control.scala 2808:40]
  wire [10:0] _GEN_140 = {{9'd0}, stride}; // @[control.scala 2809:93]
  wire [10:0] _bram_read_addr_singal_T_1 = bram_read_addr_singal + _GEN_140; // @[control.scala 2809:93]
  wire [10:0] _bram_read_addr_double_T_1 = bram_read_addr_double + _GEN_140; // @[control.scala 2810:93]
  wire [11:0] _bram_read_addr_s1_T = {1'h0,bram_read_addr_singal}; // @[Cat.scala 33:92]
  wire [11:0] _bram_read_addr_s1_T_1 = {1'h1,bram_read_addr_double}; // @[Cat.scala 33:92]
  wire [11:0] bram_read_addr_s1 = row_is_singal ? _bram_read_addr_s1_T : _bram_read_addr_s1_T_1; // @[control.scala 2812:32]
  wire [1:0] kernal_valid = {io_kernal, 1'h0}; // @[control.scala 2827:32]
  wire  _ifm_data_valid_T_1 = row_cnt < conv_row_include_pad; // @[control.scala 2830:46]
  reg  line_row_valid; // @[control.scala 2834:33]
  wire [9:0] _GEN_142 = {{8'd0}, kernal_valid}; // @[control.scala 2835:32]
  wire  line_data_valid = line_row_valid & col_cnt >= _GEN_142; // @[control.scala 2837:39]
  reg  line_data_sub_zero_valid; // @[control.scala 2838:43]
  reg  line_row_sub_zero_valid; // @[control.scala 2841:42]
  reg  line_row_sub_zero_valid_delay; // @[control.scala 2843:48]
  reg  conv_valid_s1; // @[control.scala 2849:32]
  reg  conv_valid_s2_r; // @[Reg.scala 35:20]
  reg  conv_valid_s2_r_1; // @[Reg.scala 35:20]
  wire  conv_valid_s2 = conv_valid_s2_r_1 & line_row_sub_zero_valid_delay; // @[control.scala 2850:78]
  reg  conv_valid_s1_r; // @[Reg.scala 35:20]
  reg  conv_valid_s1_r_1; // @[Reg.scala 35:20]
  reg  conv_valid_s1_r_2; // @[Reg.scala 35:20]
  wire  _conv_valid_s1_T = io_kernal ? line_row_sub_zero_valid_delay : 1'h1; // @[control.scala 2851:83]
  reg  acc_read_en_r; // @[Reg.scala 35:20]
  reg  acc_read_en_r_1; // @[Reg.scala 35:20]
  reg  acc_read_en_r_2; // @[Reg.scala 35:20]
  reg  acc_read_en_r_3; // @[Reg.scala 35:20]
  reg  acc_read_en_r_4; // @[Reg.scala 35:20]
  reg  acc_read_en_r_5; // @[Reg.scala 35:20]
  reg  acc_read_en_r_6; // @[Reg.scala 35:20]
  reg  acc_write_en_r; // @[Reg.scala 35:20]
  reg  acc_write_en; // @[Reg.scala 35:20]
  reg [11:0] acc_read_addr; // @[control.scala 2858:32]
  wire [11:0] _acc_read_addr_T_1 = acc_read_addr + 12'h1; // @[control.scala 2860:75]
  reg [11:0] acc_write_addr_r; // @[Reg.scala 35:20]
  reg [11:0] acc_write_addr_r_1; // @[Reg.scala 35:20]
  reg  io_acc_curr_data_zero_REG; // @[control.scala 2867:38]
  reg  ofm_valid_skip_act_r; // @[Reg.scala 35:20]
  reg  ofm_valid_skip_act_r_1; // @[Reg.scala 35:20]
  reg  ofm_valid_skip_act_r_2; // @[Reg.scala 35:20]
  reg  ofm_valid_skip_act_r_3; // @[Reg.scala 35:20]
  reg  ofm_valid_skip_act_r_4; // @[Reg.scala 35:20]
  reg  ofm_valid_skip_act; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_1; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_2; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_3; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_4; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_5; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_6; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_7; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_8; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_9; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_10; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_11; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_12; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_13; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_14; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_15; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_16; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_17; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_18; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_19; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_20; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_21; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_22; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_23; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_24; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_25; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_26; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act_r_27; // @[Reg.scala 35:20]
  reg  ofm_valid_after_act; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act_r; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act_r_2; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act_r_3; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act_r_4; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_skip_act; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_2; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_3; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_4; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_5; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_6; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_7; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_8; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_9; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_10; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_11; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_12; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_13; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_14; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_15; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_16; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_17; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_18; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_19; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_20; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_21; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_22; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_23; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_24; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_25; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_26; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act_r_27; // @[Reg.scala 35:20]
  reg [11:0] ofm_addr_after_act; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_1; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_2; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_3; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_4; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_5; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_6; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_7; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_8; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_9; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_10; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_11; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_12; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_13; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2_r_14; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s2; // @[Reg.scala 35:20]
  reg  ofm_done_skip_act_s1; // @[control.scala 2879:39]
  wire  ofm_done_skip_act = io_s_mod ? ofm_done_skip_act_s2 : ofm_done_skip_act_s1; // @[control.scala 2880:30]
  reg  ofm_done_after_act_r; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_1; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_2; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_3; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_4; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_5; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_6; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_7; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_8; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_9; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_10; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_11; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_12; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_13; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_14; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_15; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_16; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_17; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_18; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_19; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_20; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_21; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_22; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_23; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_24; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_25; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_26; // @[Reg.scala 35:20]
  reg  ofm_done_after_act_r_27; // @[Reg.scala 35:20]
  reg  ofm_done_after_act; // @[Reg.scala 35:20]
  wire  ofm_done = io_skip_act ? ofm_done_skip_act : ofm_done_after_act; // @[control.scala 2882:20]
  reg  io_ofm_done_REG; // @[utils.scala 19:16]
  assign io_ifmbuf_bram_addr_read_s1 = bram_read_addr_s1[11:1]; // @[control.scala 2813:53]
  assign io_ifmbuf_addr_read_sel_s1 = bram_read_addr_s1[0]; // @[control.scala 2814:52]
  assign io_ifmbuf_bram_addr_read_s2_singal = bram_read_addr_singal[10:1]; // @[control.scala 2815:64]
  assign io_ifmbuf_bram_addr_read_s2_double = bram_read_addr_double[10:1]; // @[control.scala 2816:64]
  assign io_acc_read_addr = acc_read_addr; // @[control.scala 2864:22]
  assign io_acc_write_addr = acc_write_addr_r_1; // @[control.scala 2859:30 2861:20]
  assign io_acc_read_en = acc_read_en_r_6; // @[control.scala 2855:27 2856:17]
  assign io_acc_write_en = acc_write_en; // @[control.scala 2863:20]
  assign io_acc_curr_data_zero = ~io_acc_curr_data_zero_REG; // @[control.scala 2867:30]
  assign io_ofm_addr = io_skip_act ? ofm_addr_skip_act : ofm_addr_after_act; // @[control.scala 2875:23]
  assign io_ofm_valid = io_skip_act ? ofm_valid_skip_act : ofm_valid_after_act; // @[control.scala 2871:24]
  assign io_ofm_done = io_ofm_done_REG & ~ofm_done; // @[utils.scala 19:26]
  assign io_zero_pad_valid_s1 = io_zero_pad_valid_s1_REG; // @[control.scala 2785:26]
  assign io_zero_pad_valid_s2 = io_zero_pad_valid_s2_REG; // @[control.scala 2798:25]
  always @(posedge clock) begin
    if (reset) begin // @[control.scala 2766:26]
      col_cnt <= 10'h0; // @[control.scala 2766:26]
    end else if (io_shutdown | col_cnt == conv_col_minus_stride) begin // @[control.scala 2769:19]
      col_cnt <= 10'h0;
    end else begin
      col_cnt <= _col_cnt_T_3;
    end
    if (reset) begin // @[control.scala 2767:26]
      row_cnt <= 10'h0; // @[control.scala 2767:26]
    end else if (io_shutdown) begin // @[control.scala 2770:19]
      row_cnt <= 10'h0;
    end else if (_col_cnt_T) begin // @[control.scala 2770:41]
      row_cnt <= _row_cnt_T_2;
    end
    io_zero_pad_valid_s1_REG <= zero_pad_left_and_right | zero_pad_top | zero_pad_bottom_include_top |
      zero_pad_only_bottom; // @[control.scala 2784:88]
    io_zero_pad_valid_s2_REG <= {io_zero_pad_valid_s2_hi,io_zero_pad_valid_s2_lo}; // @[Cat.scala 33:92]
    if (reset) begin // @[control.scala 2800:42]
      row_is_singal_or_double <= 1'h0; // @[control.scala 2800:42]
    end else if (io_shutdown) begin // @[control.scala 2803:35]
      row_is_singal_or_double <= 1'h0;
    end else if (_col_cnt_T) begin // @[control.scala 2803:61]
      row_is_singal_or_double <= ~row_is_singal_or_double;
    end
    if (reset) begin // @[control.scala 2807:40]
      bram_read_addr_singal <= 11'h0; // @[control.scala 2807:40]
    end else if (io_shutdown) begin // @[control.scala 2809:33]
      bram_read_addr_singal <= 11'h0;
    end else if (row_is_singal) begin // @[control.scala 2809:55]
      bram_read_addr_singal <= _bram_read_addr_singal_T_1;
    end
    if (reset) begin // @[control.scala 2808:40]
      bram_read_addr_double <= 11'h0; // @[control.scala 2808:40]
    end else if (io_shutdown) begin // @[control.scala 2810:33]
      bram_read_addr_double <= 11'h0;
    end else if (row_is_double) begin // @[control.scala 2810:55]
      bram_read_addr_double <= _bram_read_addr_double_T_1;
    end
    if (reset) begin // @[control.scala 2834:33]
      line_row_valid <= 1'h0; // @[control.scala 2834:33]
    end else begin
      line_row_valid <= row_cnt >= _GEN_142 & _ifm_data_valid_T_1; // @[control.scala 2835:20]
    end
    if (reset) begin // @[control.scala 2838:43]
      line_data_sub_zero_valid <= 1'h0; // @[control.scala 2838:43]
    end else begin
      line_data_sub_zero_valid <= line_data_valid; // @[control.scala 2839:30]
    end
    if (reset) begin // @[control.scala 2841:42]
      line_row_sub_zero_valid <= 1'h0; // @[control.scala 2841:42]
    end else begin
      line_row_sub_zero_valid <= line_row_valid; // @[control.scala 2842:29]
    end
    if (reset) begin // @[control.scala 2843:48]
      line_row_sub_zero_valid_delay <= 1'h0; // @[control.scala 2843:48]
    end else begin
      line_row_sub_zero_valid_delay <= line_row_sub_zero_valid; // @[control.scala 2844:35]
    end
    if (reset) begin // @[control.scala 2849:32]
      conv_valid_s1 <= 1'h0; // @[control.scala 2849:32]
    end else begin
      conv_valid_s1 <= conv_valid_s1_r_2 & _conv_valid_s1_T; // @[control.scala 2851:19]
    end
    if (reset) begin // @[Reg.scala 35:20]
      conv_valid_s2_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      conv_valid_s2_r <= line_data_sub_zero_valid;
    end
    if (reset) begin // @[Reg.scala 35:20]
      conv_valid_s2_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      conv_valid_s2_r_1 <= conv_valid_s2_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      conv_valid_s1_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      conv_valid_s1_r <= line_data_sub_zero_valid;
    end
    if (reset) begin // @[Reg.scala 35:20]
      conv_valid_s1_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      conv_valid_s1_r_1 <= conv_valid_s1_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      conv_valid_s1_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      conv_valid_s1_r_2 <= conv_valid_s1_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_s_mod) begin // @[control.scala 2853:22]
      acc_read_en_r <= conv_valid_s2;
    end else begin
      acc_read_en_r <= conv_valid_s1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_1 <= acc_read_en_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_2 <= acc_read_en_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_3 <= acc_read_en_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_4 <= acc_read_en_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_5 <= acc_read_en_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_read_en_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_read_en_r_6 <= acc_read_en_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_write_en_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_write_en_r <= acc_read_en_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_write_en <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      acc_write_en <= acc_write_en_r;
    end
    if (reset) begin // @[control.scala 2858:32]
      acc_read_addr <= 12'h0; // @[control.scala 2858:32]
    end else if (io_shutdown) begin // @[control.scala 2860:25]
      acc_read_addr <= 12'h0;
    end else if (acc_read_en_r_6) begin // @[control.scala 2860:47]
      acc_read_addr <= _acc_read_addr_T_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_write_addr_r <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      acc_write_addr_r <= acc_read_addr;
    end
    if (reset) begin // @[Reg.scala 35:20]
      acc_write_addr_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      acc_write_addr_r_1 <= acc_write_addr_r;
    end
    io_acc_curr_data_zero_REG <= acc_read_en_r_6; // @[control.scala 2855:27 2856:17]
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act_r <= acc_write_en;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act_r_1 <= ofm_valid_skip_act_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act_r_2 <= ofm_valid_skip_act_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act_r_3 <= ofm_valid_skip_act_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act_r_4 <= ofm_valid_skip_act_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_skip_act <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_skip_act <= ofm_valid_skip_act_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r <= ofm_valid_skip_act;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_1 <= ofm_valid_after_act_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_2 <= ofm_valid_after_act_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_3 <= ofm_valid_after_act_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_4 <= ofm_valid_after_act_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_5 <= ofm_valid_after_act_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_6 <= ofm_valid_after_act_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_7 <= ofm_valid_after_act_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_8 <= ofm_valid_after_act_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_9 <= ofm_valid_after_act_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_10 <= ofm_valid_after_act_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_11 <= ofm_valid_after_act_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_12 <= ofm_valid_after_act_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_13 <= ofm_valid_after_act_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_14 <= ofm_valid_after_act_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_15 <= ofm_valid_after_act_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_16 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_16 <= ofm_valid_after_act_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_17 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_17 <= ofm_valid_after_act_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_18 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_18 <= ofm_valid_after_act_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_19 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_19 <= ofm_valid_after_act_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_20 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_20 <= ofm_valid_after_act_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_21 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_21 <= ofm_valid_after_act_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_22 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_22 <= ofm_valid_after_act_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_23 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_23 <= ofm_valid_after_act_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_24 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_24 <= ofm_valid_after_act_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_25 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_25 <= ofm_valid_after_act_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_26 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_26 <= ofm_valid_after_act_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act_r_27 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act_r_27 <= ofm_valid_after_act_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_valid_after_act <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_valid_after_act <= ofm_valid_after_act_r_27;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act_r <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act_r <= acc_write_addr_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act_r_1 <= ofm_addr_skip_act_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act_r_2 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act_r_2 <= ofm_addr_skip_act_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act_r_3 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act_r_3 <= ofm_addr_skip_act_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act_r_4 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act_r_4 <= ofm_addr_skip_act_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_skip_act <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_skip_act <= ofm_addr_skip_act_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r <= ofm_addr_skip_act;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_1 <= ofm_addr_after_act_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_2 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_2 <= ofm_addr_after_act_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_3 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_3 <= ofm_addr_after_act_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_4 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_4 <= ofm_addr_after_act_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_5 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_5 <= ofm_addr_after_act_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_6 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_6 <= ofm_addr_after_act_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_7 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_7 <= ofm_addr_after_act_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_8 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_8 <= ofm_addr_after_act_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_9 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_9 <= ofm_addr_after_act_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_10 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_10 <= ofm_addr_after_act_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_11 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_11 <= ofm_addr_after_act_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_12 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_12 <= ofm_addr_after_act_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_13 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_13 <= ofm_addr_after_act_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_14 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_14 <= ofm_addr_after_act_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_15 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_15 <= ofm_addr_after_act_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_16 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_16 <= ofm_addr_after_act_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_17 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_17 <= ofm_addr_after_act_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_18 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_18 <= ofm_addr_after_act_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_19 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_19 <= ofm_addr_after_act_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_20 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_20 <= ofm_addr_after_act_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_21 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_21 <= ofm_addr_after_act_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_22 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_22 <= ofm_addr_after_act_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_23 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_23 <= ofm_addr_after_act_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_24 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_24 <= ofm_addr_after_act_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_25 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_25 <= ofm_addr_after_act_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_26 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_26 <= ofm_addr_after_act_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act_r_27 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act_r_27 <= ofm_addr_after_act_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_addr_after_act <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_addr_after_act <= ofm_addr_after_act_r_27;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r <= line_row_sub_zero_valid;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_1 <= ofm_done_skip_act_s2_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_2 <= ofm_done_skip_act_s2_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_3 <= ofm_done_skip_act_s2_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_4 <= ofm_done_skip_act_s2_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_5 <= ofm_done_skip_act_s2_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_6 <= ofm_done_skip_act_s2_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_7 <= ofm_done_skip_act_s2_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_8 <= ofm_done_skip_act_s2_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_9 <= ofm_done_skip_act_s2_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_10 <= ofm_done_skip_act_s2_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_11 <= ofm_done_skip_act_s2_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_12 <= ofm_done_skip_act_s2_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_13 <= ofm_done_skip_act_s2_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2_r_14 <= ofm_done_skip_act_s2_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_skip_act_s2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_skip_act_s2 <= ofm_done_skip_act_s2_r_14;
    end
    ofm_done_skip_act_s1 <= ofm_done_skip_act_s2; // @[control.scala 2879:39]
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_s_mod) begin // @[control.scala 2880:30]
      ofm_done_after_act_r <= ofm_done_skip_act_s2;
    end else begin
      ofm_done_after_act_r <= ofm_done_skip_act_s1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_1 <= ofm_done_after_act_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_2 <= ofm_done_after_act_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_3 <= ofm_done_after_act_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_4 <= ofm_done_after_act_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_5 <= ofm_done_after_act_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_6 <= ofm_done_after_act_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_7 <= ofm_done_after_act_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_8 <= ofm_done_after_act_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_9 <= ofm_done_after_act_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_10 <= ofm_done_after_act_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_11 <= ofm_done_after_act_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_12 <= ofm_done_after_act_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_13 <= ofm_done_after_act_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_14 <= ofm_done_after_act_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_15 <= ofm_done_after_act_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_16 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_16 <= ofm_done_after_act_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_17 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_17 <= ofm_done_after_act_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_18 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_18 <= ofm_done_after_act_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_19 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_19 <= ofm_done_after_act_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_20 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_20 <= ofm_done_after_act_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_21 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_21 <= ofm_done_after_act_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_22 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_22 <= ofm_done_after_act_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_23 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_23 <= ofm_done_after_act_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_24 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_24 <= ofm_done_after_act_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_25 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_25 <= ofm_done_after_act_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_26 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_26 <= ofm_done_after_act_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act_r_27 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act_r_27 <= ofm_done_after_act_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_done_after_act <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_done_after_act <= ofm_done_after_act_r_27;
    end
    if (reset) begin // @[utils.scala 19:16]
      io_ofm_done_REG <= 1'h0; // @[utils.scala 19:16]
    end else if (io_skip_act) begin // @[control.scala 2882:20]
      if (io_s_mod) begin // @[control.scala 2880:30]
        io_ofm_done_REG <= ofm_done_skip_act_s2;
      end else begin
        io_ofm_done_REG <= ofm_done_skip_act_s1;
      end
    end else begin
      io_ofm_done_REG <= ofm_done_after_act;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  col_cnt = _RAND_0[9:0];
  _RAND_1 = {1{`RANDOM}};
  row_cnt = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  io_zero_pad_valid_s1_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_zero_pad_valid_s2_REG = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  row_is_singal_or_double = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  bram_read_addr_singal = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  bram_read_addr_double = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  line_row_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  line_data_sub_zero_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  line_row_sub_zero_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  line_row_sub_zero_valid_delay = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  conv_valid_s1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  conv_valid_s2_r = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  conv_valid_s2_r_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  conv_valid_s1_r = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  conv_valid_s1_r_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  conv_valid_s1_r_2 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  acc_read_en_r = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  acc_read_en_r_1 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  acc_read_en_r_2 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  acc_read_en_r_3 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  acc_read_en_r_4 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  acc_read_en_r_5 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  acc_read_en_r_6 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  acc_write_en_r = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  acc_write_en = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  acc_read_addr = _RAND_26[11:0];
  _RAND_27 = {1{`RANDOM}};
  acc_write_addr_r = _RAND_27[11:0];
  _RAND_28 = {1{`RANDOM}};
  acc_write_addr_r_1 = _RAND_28[11:0];
  _RAND_29 = {1{`RANDOM}};
  io_acc_curr_data_zero_REG = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  ofm_valid_skip_act_r = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  ofm_valid_skip_act_r_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  ofm_valid_skip_act_r_2 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  ofm_valid_skip_act_r_3 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  ofm_valid_skip_act_r_4 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ofm_valid_skip_act = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  ofm_valid_after_act_r = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ofm_valid_after_act_r_1 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ofm_valid_after_act_r_2 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  ofm_valid_after_act_r_3 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  ofm_valid_after_act_r_4 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ofm_valid_after_act_r_5 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  ofm_valid_after_act_r_6 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  ofm_valid_after_act_r_7 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  ofm_valid_after_act_r_8 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  ofm_valid_after_act_r_9 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ofm_valid_after_act_r_10 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ofm_valid_after_act_r_11 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  ofm_valid_after_act_r_12 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ofm_valid_after_act_r_13 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ofm_valid_after_act_r_14 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ofm_valid_after_act_r_15 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ofm_valid_after_act_r_16 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ofm_valid_after_act_r_17 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ofm_valid_after_act_r_18 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ofm_valid_after_act_r_19 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ofm_valid_after_act_r_20 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  ofm_valid_after_act_r_21 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  ofm_valid_after_act_r_22 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  ofm_valid_after_act_r_23 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  ofm_valid_after_act_r_24 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  ofm_valid_after_act_r_25 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  ofm_valid_after_act_r_26 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  ofm_valid_after_act_r_27 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  ofm_valid_after_act = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  ofm_addr_skip_act_r = _RAND_65[11:0];
  _RAND_66 = {1{`RANDOM}};
  ofm_addr_skip_act_r_1 = _RAND_66[11:0];
  _RAND_67 = {1{`RANDOM}};
  ofm_addr_skip_act_r_2 = _RAND_67[11:0];
  _RAND_68 = {1{`RANDOM}};
  ofm_addr_skip_act_r_3 = _RAND_68[11:0];
  _RAND_69 = {1{`RANDOM}};
  ofm_addr_skip_act_r_4 = _RAND_69[11:0];
  _RAND_70 = {1{`RANDOM}};
  ofm_addr_skip_act = _RAND_70[11:0];
  _RAND_71 = {1{`RANDOM}};
  ofm_addr_after_act_r = _RAND_71[11:0];
  _RAND_72 = {1{`RANDOM}};
  ofm_addr_after_act_r_1 = _RAND_72[11:0];
  _RAND_73 = {1{`RANDOM}};
  ofm_addr_after_act_r_2 = _RAND_73[11:0];
  _RAND_74 = {1{`RANDOM}};
  ofm_addr_after_act_r_3 = _RAND_74[11:0];
  _RAND_75 = {1{`RANDOM}};
  ofm_addr_after_act_r_4 = _RAND_75[11:0];
  _RAND_76 = {1{`RANDOM}};
  ofm_addr_after_act_r_5 = _RAND_76[11:0];
  _RAND_77 = {1{`RANDOM}};
  ofm_addr_after_act_r_6 = _RAND_77[11:0];
  _RAND_78 = {1{`RANDOM}};
  ofm_addr_after_act_r_7 = _RAND_78[11:0];
  _RAND_79 = {1{`RANDOM}};
  ofm_addr_after_act_r_8 = _RAND_79[11:0];
  _RAND_80 = {1{`RANDOM}};
  ofm_addr_after_act_r_9 = _RAND_80[11:0];
  _RAND_81 = {1{`RANDOM}};
  ofm_addr_after_act_r_10 = _RAND_81[11:0];
  _RAND_82 = {1{`RANDOM}};
  ofm_addr_after_act_r_11 = _RAND_82[11:0];
  _RAND_83 = {1{`RANDOM}};
  ofm_addr_after_act_r_12 = _RAND_83[11:0];
  _RAND_84 = {1{`RANDOM}};
  ofm_addr_after_act_r_13 = _RAND_84[11:0];
  _RAND_85 = {1{`RANDOM}};
  ofm_addr_after_act_r_14 = _RAND_85[11:0];
  _RAND_86 = {1{`RANDOM}};
  ofm_addr_after_act_r_15 = _RAND_86[11:0];
  _RAND_87 = {1{`RANDOM}};
  ofm_addr_after_act_r_16 = _RAND_87[11:0];
  _RAND_88 = {1{`RANDOM}};
  ofm_addr_after_act_r_17 = _RAND_88[11:0];
  _RAND_89 = {1{`RANDOM}};
  ofm_addr_after_act_r_18 = _RAND_89[11:0];
  _RAND_90 = {1{`RANDOM}};
  ofm_addr_after_act_r_19 = _RAND_90[11:0];
  _RAND_91 = {1{`RANDOM}};
  ofm_addr_after_act_r_20 = _RAND_91[11:0];
  _RAND_92 = {1{`RANDOM}};
  ofm_addr_after_act_r_21 = _RAND_92[11:0];
  _RAND_93 = {1{`RANDOM}};
  ofm_addr_after_act_r_22 = _RAND_93[11:0];
  _RAND_94 = {1{`RANDOM}};
  ofm_addr_after_act_r_23 = _RAND_94[11:0];
  _RAND_95 = {1{`RANDOM}};
  ofm_addr_after_act_r_24 = _RAND_95[11:0];
  _RAND_96 = {1{`RANDOM}};
  ofm_addr_after_act_r_25 = _RAND_96[11:0];
  _RAND_97 = {1{`RANDOM}};
  ofm_addr_after_act_r_26 = _RAND_97[11:0];
  _RAND_98 = {1{`RANDOM}};
  ofm_addr_after_act_r_27 = _RAND_98[11:0];
  _RAND_99 = {1{`RANDOM}};
  ofm_addr_after_act = _RAND_99[11:0];
  _RAND_100 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_1 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_2 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_3 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_4 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_5 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_6 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_7 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_8 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_9 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_10 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_11 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_12 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_13 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  ofm_done_skip_act_s2_r_14 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  ofm_done_skip_act_s2 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  ofm_done_skip_act_s1 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  ofm_done_after_act_r = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  ofm_done_after_act_r_1 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  ofm_done_after_act_r_2 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  ofm_done_after_act_r_3 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  ofm_done_after_act_r_4 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  ofm_done_after_act_r_5 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  ofm_done_after_act_r_6 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  ofm_done_after_act_r_7 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  ofm_done_after_act_r_8 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  ofm_done_after_act_r_9 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  ofm_done_after_act_r_10 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  ofm_done_after_act_r_11 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  ofm_done_after_act_r_12 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  ofm_done_after_act_r_13 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  ofm_done_after_act_r_14 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  ofm_done_after_act_r_15 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  ofm_done_after_act_r_16 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  ofm_done_after_act_r_17 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  ofm_done_after_act_r_18 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  ofm_done_after_act_r_19 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  ofm_done_after_act_r_20 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  ofm_done_after_act_r_21 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  ofm_done_after_act_r_22 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  ofm_done_after_act_r_23 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  ofm_done_after_act_r_24 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  ofm_done_after_act_r_25 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  ofm_done_after_act_r_26 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  ofm_done_after_act_r_27 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  ofm_done_after_act = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  io_ofm_done_REG = _RAND_146[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DMA_Master(
  input         clock,
  input         reset,
  input         io_send_enable,
  output        io_send_done,
  input  [31:0] io_dma_addr,
  input  [15:0] io_dma_len,
  output        io_dma_wvalid,
  input         io_dma_wbusy,
  input         io_dma_wready,
  output        io_dma_wareq,
  output [31:0] io_dma_waddr,
  output [15:0] io_dma_wsize,
  output [63:0] io_dma_wdata,
  input  [16:0] io_addr_start,
  input  [16:0] io_addr_end,
  output [16:0] io_read_addr,
  input  [63:0] io_read_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [16:0] addr; // @[DMA_Master_and_slave.scala 35:23]
  reg  last_d; // @[DMA_Master_and_slave.scala 38:25]
  reg  send_enable_flag; // @[DMA_Master_and_slave.scala 45:35]
  reg  send_enable_u_REG; // @[utils.scala 10:17]
  wire  send_enable_u = ~send_enable_u_REG & io_send_enable; // @[utils.scala 10:27]
  reg  dma_wareq; // @[DMA_Master_and_slave.scala 68:28]
  wire  _dma_wareq_T_5 = dma_wareq & io_dma_wbusy ? 1'h0 : dma_wareq; // @[DMA_Master_and_slave.scala 70:75]
  reg [8:0] addr_cnt; // @[DMA_Master_and_slave.scala 71:27]
  wire [8:0] _addr_cnt_T_3 = addr_cnt + 9'h1; // @[DMA_Master_and_slave.scala 72:103]
  wire [16:0] _last_T_1 = io_addr_end - io_addr_start; // @[DMA_Master_and_slave.scala 82:40]
  wire [16:0] _last_T_3 = _last_T_1 - 17'h1; // @[DMA_Master_and_slave.scala 82:56]
  wire  last = addr == _last_T_3; // @[DMA_Master_and_slave.scala 82:23]
  wire [16:0] _addr_T_1 = addr + 17'h1; // @[DMA_Master_and_slave.scala 84:50]
  wire  addr_en = addr_cnt > 9'h3 & addr_cnt < 9'h104; // @[DMA_Master_and_slave.scala 86:33]
  reg  r_dma_wvalid; // @[DMA_Master_and_slave.scala 87:31]
  assign io_send_done = last_d; // @[DMA_Master_and_slave.scala 39:25 40:15]
  assign io_dma_wvalid = r_dma_wvalid; // @[DMA_Master_and_slave.scala 89:19]
  assign io_dma_wareq = dma_wareq; // @[DMA_Master_and_slave.scala 69:18]
  assign io_dma_waddr = io_dma_addr; // @[DMA_Master_and_slave.scala 33:18]
  assign io_dma_wsize = io_dma_len; // @[DMA_Master_and_slave.scala 32:18]
  assign io_dma_wdata = io_read_data; // @[DMA_Master_and_slave.scala 83:22]
  assign io_read_addr = addr + io_addr_start; // @[DMA_Master_and_slave.scala 49:26]
  always @(posedge clock) begin
    if (reset) begin // @[DMA_Master_and_slave.scala 35:23]
      addr <= 17'h0; // @[DMA_Master_and_slave.scala 35:23]
    end else if (last) begin // @[DMA_Master_and_slave.scala 84:20]
      addr <= 17'h0;
    end else if (addr_en) begin // @[DMA_Master_and_slave.scala 84:35]
      addr <= _addr_T_1;
    end
    last_d <= addr == _last_T_3; // @[DMA_Master_and_slave.scala 82:23]
    if (reset) begin // @[DMA_Master_and_slave.scala 45:35]
      send_enable_flag <= 1'h0; // @[DMA_Master_and_slave.scala 45:35]
    end else if (io_dma_wareq) begin // @[DMA_Master_and_slave.scala 46:28]
      send_enable_flag <= 1'h0;
    end else begin
      send_enable_flag <= send_enable_u | send_enable_flag;
    end
    if (reset) begin // @[utils.scala 10:17]
      send_enable_u_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      send_enable_u_REG <= io_send_enable; // @[utils.scala 10:17]
    end
    if (reset) begin // @[DMA_Master_and_slave.scala 68:28]
      dma_wareq <= 1'h0; // @[DMA_Master_and_slave.scala 68:28]
    end else begin
      dma_wareq <= send_enable_flag & ~io_dma_wbusy | _dma_wareq_T_5; // @[DMA_Master_and_slave.scala 70:15]
    end
    if (reset) begin // @[DMA_Master_and_slave.scala 71:27]
      addr_cnt <= 9'h0; // @[DMA_Master_and_slave.scala 71:27]
    end else if (last) begin // @[DMA_Master_and_slave.scala 72:20]
      addr_cnt <= 9'h0;
    end else if (io_dma_wbusy & io_dma_wready) begin // @[DMA_Master_and_slave.scala 72:35]
      if (addr_cnt == 9'h108) begin // @[DMA_Master_and_slave.scala 72:68]
        addr_cnt <= 9'h4;
      end else begin
        addr_cnt <= _addr_cnt_T_3;
      end
    end else begin
      addr_cnt <= 9'h0;
    end
    if (reset) begin // @[DMA_Master_and_slave.scala 87:31]
      r_dma_wvalid <= 1'h0; // @[DMA_Master_and_slave.scala 87:31]
    end else begin
      r_dma_wvalid <= addr_en; // @[DMA_Master_and_slave.scala 88:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[16:0];
  _RAND_1 = {1{`RANDOM}};
  last_d = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  send_enable_flag = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  send_enable_u_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  dma_wareq = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  addr_cnt = _RAND_5[8:0];
  _RAND_6 = {1{`RANDOM}};
  r_dma_wvalid = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DMA_Slave(
  input         clock,
  input         reset,
  input         io_recv_enable,
  output        io_recv_done,
  input  [31:0] io_dma_addr,
  input  [15:0] io_dma_len,
  input         io_dma_rvalid,
  input         io_dma_rbusy,
  output        io_dma_rareq,
  output [31:0] io_dma_raddr,
  output [15:0] io_dma_rsize,
  input  [63:0] io_dma_rdata,
  output [63:0] io_write_data,
  output        io_write_enable
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  dma_rbusy_downedge_REG; // @[utils.scala 19:16]
  wire  _dma_rbusy_downedge_T = ~io_dma_rbusy; // @[utils.scala 19:29]
  wire  dma_rbusy_downedge = dma_rbusy_downedge_REG & ~io_dma_rbusy; // @[utils.scala 19:26]
  wire  clr = reset | dma_rbusy_downedge; // @[DMA_Master_and_slave.scala 124:27]
  wire  write_enable = io_dma_rbusy & io_dma_rvalid; // @[DMA_Master_and_slave.scala 127:37]
  reg [63:0] r_write_data; // @[DMA_Master_and_slave.scala 132:35]
  reg  r_write_enable; // @[DMA_Master_and_slave.scala 133:37]
  reg  recv_enable_up_REG; // @[utils.scala 10:17]
  wire  recv_enable_up = ~recv_enable_up_REG & io_recv_enable; // @[utils.scala 10:27]
  reg  recv_enable_flag; // @[DMA_Master_and_slave.scala 137:39]
  reg  dma_rareq; // @[DMA_Master_and_slave.scala 139:32]
  wire  _dma_rareq_T_3 = io_dma_rareq & io_dma_rbusy ? 1'h0 : io_dma_rareq; // @[DMA_Master_and_slave.scala 140:71]
  assign io_recv_done = dma_rbusy_downedge_REG & ~io_dma_rbusy; // @[utils.scala 19:26]
  assign io_dma_rareq = dma_rareq; // @[DMA_Master_and_slave.scala 143:22]
  assign io_dma_raddr = io_dma_addr; // @[DMA_Master_and_slave.scala 116:18]
  assign io_dma_rsize = io_dma_len; // @[DMA_Master_and_slave.scala 117:18]
  assign io_write_data = r_write_data; // @[DMA_Master_and_slave.scala 160:27]
  assign io_write_enable = r_write_enable; // @[DMA_Master_and_slave.scala 161:28]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 19:16]
      dma_rbusy_downedge_REG <= 1'h0; // @[utils.scala 19:16]
    end else begin
      dma_rbusy_downedge_REG <= io_dma_rbusy; // @[utils.scala 19:16]
    end
    if (clr) begin // @[DMA_Master_and_slave.scala 132:35]
      r_write_data <= 64'h0; // @[DMA_Master_and_slave.scala 132:35]
    end else begin
      r_write_data <= io_dma_rdata; // @[DMA_Master_and_slave.scala 158:26]
    end
    if (clr) begin // @[DMA_Master_and_slave.scala 133:37]
      r_write_enable <= 1'h0; // @[DMA_Master_and_slave.scala 133:37]
    end else begin
      r_write_enable <= write_enable; // @[DMA_Master_and_slave.scala 159:28]
    end
    if (clr) begin // @[utils.scala 10:17]
      recv_enable_up_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      recv_enable_up_REG <= io_recv_enable; // @[utils.scala 10:17]
    end
    if (clr) begin // @[DMA_Master_and_slave.scala 137:39]
      recv_enable_flag <= 1'h0; // @[DMA_Master_and_slave.scala 137:39]
    end else if (io_dma_rareq) begin // @[DMA_Master_and_slave.scala 138:32]
      recv_enable_flag <= 1'h0;
    end else begin
      recv_enable_flag <= recv_enable_up | recv_enable_flag;
    end
    if (clr) begin // @[DMA_Master_and_slave.scala 139:32]
      dma_rareq <= 1'h0; // @[DMA_Master_and_slave.scala 139:32]
    end else begin
      dma_rareq <= recv_enable_flag & _dma_rbusy_downedge_T | _dma_rareq_T_3; // @[DMA_Master_and_slave.scala 140:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dma_rbusy_downedge_REG = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  r_write_data = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  r_write_enable = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  recv_enable_up_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  recv_enable_flag = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  dma_rareq = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ctrl_task_state(
  input   clock,
  input   reset,
  input   io_start_signal,
  input   io_done_signal,
  output  io_running
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] curr_state; // @[control.scala 3010:29]
  reg  running_state; // @[control.scala 3033:32]
  assign io_running = running_state; // @[control.scala 3035:16]
  always @(posedge clock) begin
    if (reset) begin // @[control.scala 3010:29]
      curr_state <= 2'h0; // @[control.scala 3010:29]
    end else if (2'h0 == curr_state) begin // @[control.scala 3013:24]
      if (io_start_signal) begin // @[control.scala 3015:35]
        curr_state <= 2'h1; // @[control.scala 3016:28]
      end else begin
        curr_state <= 2'h0; // @[control.scala 3018:28]
      end
    end else if (2'h1 == curr_state) begin // @[control.scala 3013:24]
      if (io_done_signal) begin // @[control.scala 3022:34]
        curr_state <= 2'h2; // @[control.scala 3023:28]
      end else begin
        curr_state <= 2'h1; // @[control.scala 3025:28]
      end
    end else if (2'h2 == curr_state) begin // @[control.scala 3013:24]
      curr_state <= 2'h0; // @[control.scala 3029:24]
    end
    if (reset) begin // @[control.scala 3033:32]
      running_state <= 1'h0; // @[control.scala 3033:32]
    end else begin
      running_state <= curr_state == 2'h1; // @[control.scala 3034:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  running_state = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ctrl_task_state_1(
  input   clock,
  input   reset,
  input   io_start_signal,
  input   io_done_signal,
  output  io_running
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] curr_state; // @[control.scala 3010:29]
  reg  running_state; // @[control.scala 3033:32]
  wire  _running_state_T_3 = curr_state == 2'h1 ? 1'h0 : 1'h1; // @[control.scala 3034:25]
  assign io_running = running_state; // @[control.scala 3035:16]
  always @(posedge clock) begin
    if (reset) begin // @[control.scala 3010:29]
      curr_state <= 2'h0; // @[control.scala 3010:29]
    end else if (2'h0 == curr_state) begin // @[control.scala 3013:24]
      if (io_start_signal) begin // @[control.scala 3015:35]
        curr_state <= 2'h1; // @[control.scala 3016:28]
      end else begin
        curr_state <= 2'h0; // @[control.scala 3018:28]
      end
    end else if (2'h1 == curr_state) begin // @[control.scala 3013:24]
      if (io_done_signal) begin // @[control.scala 3022:34]
        curr_state <= 2'h2; // @[control.scala 3023:28]
      end else begin
        curr_state <= 2'h1; // @[control.scala 3025:28]
      end
    end else if (2'h2 == curr_state) begin // @[control.scala 3013:24]
      curr_state <= 2'h0; // @[control.scala 3029:24]
    end
    running_state <= reset | _running_state_T_3; // @[control.scala 3033:{32,32} 3034:19]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  curr_state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  running_state = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module generate_ctrl_signal(
  input   clock,
  input   reset,
  input   io_recv_enable,
  input   io_send_enable,
  input   io_conv_start,
  input   io_bottleneck_add_enable,
  input   io_recv_done,
  input   io_send_done,
  input   io_conv_done,
  input   io_bottleneck_add_done,
  output  io_conv_shutdown,
  output  io_bn_add_working,
  input   io_task_valid,
  output  io_ap_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_task_state_recv_clock; // @[control.scala 2984:38]
  wire  ctrl_task_state_recv_reset; // @[control.scala 2984:38]
  wire  ctrl_task_state_recv_io_start_signal; // @[control.scala 2984:38]
  wire  ctrl_task_state_recv_io_done_signal; // @[control.scala 2984:38]
  wire  ctrl_task_state_recv_io_running; // @[control.scala 2984:38]
  wire  ctrl_task_state_conv_clock; // @[control.scala 2988:38]
  wire  ctrl_task_state_conv_reset; // @[control.scala 2988:38]
  wire  ctrl_task_state_conv_io_start_signal; // @[control.scala 2988:38]
  wire  ctrl_task_state_conv_io_done_signal; // @[control.scala 2988:38]
  wire  ctrl_task_state_conv_io_running; // @[control.scala 2988:38]
  wire  ctrl_task_state_send_clock; // @[control.scala 2992:38]
  wire  ctrl_task_state_send_reset; // @[control.scala 2992:38]
  wire  ctrl_task_state_send_io_start_signal; // @[control.scala 2992:38]
  wire  ctrl_task_state_send_io_done_signal; // @[control.scala 2992:38]
  wire  ctrl_task_state_send_io_running; // @[control.scala 2992:38]
  wire  ctrl_task_state_bn_clock; // @[control.scala 2996:36]
  wire  ctrl_task_state_bn_reset; // @[control.scala 2996:36]
  wire  ctrl_task_state_bn_io_start_signal; // @[control.scala 2996:36]
  wire  ctrl_task_state_bn_io_done_signal; // @[control.scala 2996:36]
  wire  ctrl_task_state_bn_io_running; // @[control.scala 2996:36]
  reg [3:0] task_reg; // @[control.scala 2972:27]
  wire [3:0] task_ctrl_line = {io_recv_enable,io_send_enable,io_conv_start,io_bottleneck_add_enable}; // @[Cat.scala 33:92]
  wire  _task_done_T = task_reg == 4'h8; // @[control.scala 2977:51]
  wire  _task_done_T_1 = task_reg == 4'h4; // @[control.scala 2977:93]
  wire  _task_done_T_2 = task_reg == 4'h2; // @[control.scala 2977:135]
  wire  _task_done_T_3 = task_reg == 4'ha; // @[control.scala 2977:177]
  wire  _task_done_T_4 = task_reg == 4'h9; // @[control.scala 2977:219]
  wire  _task_done_T_5 = task_reg == 4'h1; // @[control.scala 2977:261]
  wire  _task_done_T_7 = _task_done_T_4 ? io_recv_done : _task_done_T_5 & io_bottleneck_add_done; // @[Mux.scala 101:16]
  wire  _task_done_T_8 = _task_done_T_3 ? io_recv_done : _task_done_T_7; // @[Mux.scala 101:16]
  wire  _task_done_T_9 = _task_done_T_2 ? io_conv_done : _task_done_T_8; // @[Mux.scala 101:16]
  wire  _task_done_T_10 = _task_done_T_1 ? io_send_done : _task_done_T_9; // @[Mux.scala 101:16]
  wire  task_done = _task_done_T ? io_recv_done : _task_done_T_10; // @[Mux.scala 101:16]
  reg  ap_done_reg; // @[control.scala 2979:30]
  ctrl_task_state ctrl_task_state_recv ( // @[control.scala 2984:38]
    .clock(ctrl_task_state_recv_clock),
    .reset(ctrl_task_state_recv_reset),
    .io_start_signal(ctrl_task_state_recv_io_start_signal),
    .io_done_signal(ctrl_task_state_recv_io_done_signal),
    .io_running(ctrl_task_state_recv_io_running)
  );
  ctrl_task_state_1 ctrl_task_state_conv ( // @[control.scala 2988:38]
    .clock(ctrl_task_state_conv_clock),
    .reset(ctrl_task_state_conv_reset),
    .io_start_signal(ctrl_task_state_conv_io_start_signal),
    .io_done_signal(ctrl_task_state_conv_io_done_signal),
    .io_running(ctrl_task_state_conv_io_running)
  );
  ctrl_task_state ctrl_task_state_send ( // @[control.scala 2992:38]
    .clock(ctrl_task_state_send_clock),
    .reset(ctrl_task_state_send_reset),
    .io_start_signal(ctrl_task_state_send_io_start_signal),
    .io_done_signal(ctrl_task_state_send_io_done_signal),
    .io_running(ctrl_task_state_send_io_running)
  );
  ctrl_task_state ctrl_task_state_bn ( // @[control.scala 2996:36]
    .clock(ctrl_task_state_bn_clock),
    .reset(ctrl_task_state_bn_reset),
    .io_start_signal(ctrl_task_state_bn_io_start_signal),
    .io_done_signal(ctrl_task_state_bn_io_done_signal),
    .io_running(ctrl_task_state_bn_io_running)
  );
  assign io_conv_shutdown = ctrl_task_state_conv_io_running; // @[control.scala 2991:22]
  assign io_bn_add_working = ctrl_task_state_bn_io_running; // @[control.scala 2999:23]
  assign io_ap_done = ap_done_reg; // @[control.scala 2980:16]
  assign ctrl_task_state_recv_clock = clock;
  assign ctrl_task_state_recv_reset = reset;
  assign ctrl_task_state_recv_io_start_signal = io_recv_enable; // @[control.scala 2985:42]
  assign ctrl_task_state_recv_io_done_signal = io_recv_done; // @[control.scala 2986:41]
  assign ctrl_task_state_conv_clock = clock;
  assign ctrl_task_state_conv_reset = reset;
  assign ctrl_task_state_conv_io_start_signal = io_conv_start; // @[control.scala 2989:42]
  assign ctrl_task_state_conv_io_done_signal = io_conv_done; // @[control.scala 2990:41]
  assign ctrl_task_state_send_clock = clock;
  assign ctrl_task_state_send_reset = reset;
  assign ctrl_task_state_send_io_start_signal = io_send_enable; // @[control.scala 2993:42]
  assign ctrl_task_state_send_io_done_signal = io_send_done; // @[control.scala 2994:41]
  assign ctrl_task_state_bn_clock = clock;
  assign ctrl_task_state_bn_reset = reset;
  assign ctrl_task_state_bn_io_start_signal = io_bottleneck_add_enable; // @[control.scala 2997:40]
  assign ctrl_task_state_bn_io_done_signal = io_bottleneck_add_done; // @[control.scala 2998:39]
  always @(posedge clock) begin
    if (reset) begin // @[control.scala 2972:27]
      task_reg <= 4'h0; // @[control.scala 2972:27]
    end else if (io_task_valid) begin // @[control.scala 2974:20]
      task_reg <= task_ctrl_line;
    end
    if (reset) begin // @[control.scala 2979:30]
      ap_done_reg <= 1'h0; // @[control.scala 2979:30]
    end else if (io_task_valid) begin // @[control.scala 2981:23]
      ap_done_reg <= 1'h0;
    end else begin
      ap_done_reg <= task_done | ap_done_reg;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  task_reg = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  ap_done_reg = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axis_buf_sel(
  input  [1:0]  io_axis_buf_sel,
  input  [63:0] io_write_data,
  input         io_write_enable,
  output [63:0] io_write_data_ifm,
  output        io_write_enable_ifm,
  output [63:0] io_write_data_weight,
  output        io_write_enable_weight,
  output [63:0] io_write_data_bias,
  output        io_write_enable_bias
);
  wire  sel_ifm = io_axis_buf_sel == 2'h0; // @[DMA_Master_and_slave.scala 196:32]
  wire  sel_weight = io_axis_buf_sel == 2'h1; // @[DMA_Master_and_slave.scala 197:35]
  wire  sel_bias = io_axis_buf_sel == 2'h2; // @[DMA_Master_and_slave.scala 198:33]
  assign io_write_data_ifm = sel_ifm ? io_write_data : 64'h0; // @[DMA_Master_and_slave.scala 202:29]
  assign io_write_enable_ifm = sel_ifm & io_write_enable; // @[DMA_Master_and_slave.scala 203:31]
  assign io_write_data_weight = sel_weight ? io_write_data : 64'h0; // @[DMA_Master_and_slave.scala 206:32]
  assign io_write_enable_weight = sel_weight & io_write_enable; // @[DMA_Master_and_slave.scala 207:34]
  assign io_write_data_bias = sel_bias ? io_write_data : 64'h0; // @[DMA_Master_and_slave.scala 210:30]
  assign io_write_enable_bias = sel_bias & io_write_enable; // @[DMA_Master_and_slave.scala 211:32]
endmodule
module TPRAM_WRAP(
  input         clock,
  input         io_wen,
  input         io_ren,
  input  [10:0] io_waddr,
  input  [10:0] io_raddr,
  input  [15:0] io_wdata,
  output [15:0] io_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  tpram_CLKA; // @[utils.scala 218:23]
  wire  tpram_CLKB; // @[utils.scala 218:23]
  wire  tpram_CENB; // @[utils.scala 218:23]
  wire  tpram_CENA; // @[utils.scala 218:23]
  wire [10:0] tpram_AB; // @[utils.scala 218:23]
  wire [10:0] tpram_AA; // @[utils.scala 218:23]
  wire [15:0] tpram_DB; // @[utils.scala 218:23]
  wire [15:0] tpram_QA; // @[utils.scala 218:23]
  reg  rd_en; // @[utils.scala 219:46]
  reg [15:0] rdata_reg; // @[Reg.scala 19:16]
  TPRAM #(.DATA_WIDTH(16), .DEPTH(2048), .RAM_STYLE_VAL("block")) tpram ( // @[utils.scala 218:23]
    .CLKA(tpram_CLKA),
    .CLKB(tpram_CLKB),
    .CENB(tpram_CENB),
    .CENA(tpram_CENA),
    .AB(tpram_AB),
    .AA(tpram_AA),
    .DB(tpram_DB),
    .QA(tpram_QA)
  );
  assign io_rdata = ~rd_en ? rdata_reg : tpram_QA; // @[utils.scala 230:12]
  assign tpram_CLKA = clock; // @[utils.scala 222:19]
  assign tpram_CLKB = clock; // @[utils.scala 223:19]
  assign tpram_CENB = ~io_wen; // @[utils.scala 224:22]
  assign tpram_CENA = ~io_ren; // @[utils.scala 225:22]
  assign tpram_AB = io_waddr; // @[utils.scala 226:17]
  assign tpram_AA = io_raddr; // @[utils.scala 227:17]
  assign tpram_DB = io_wdata; // @[utils.scala 228:17]
  always @(posedge clock) begin
    rd_en <= io_ren; // @[utils.scala 219:46]
    if (rd_en) begin // @[Reg.scala 20:18]
      rdata_reg <= tpram_QA; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_en = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rdata_reg = _RAND_1[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IfmBuffer(
  input         clock,
  input         reset,
  input  [10:0] io_ifmbuf_bram_addr_read_s1,
  input         io_ifmbuf_bram_addr_read_sel_s1,
  input  [9:0]  io_ifmbuf_bram_addr_read_s2_singal,
  input  [9:0]  io_ifmbuf_bram_addr_read_s2_double,
  input         io_bram_en_write,
  input         io_upsample_enable,
  input         io_recv_done,
  input         io_buf_sel,
  input         io_s_mod,
  input  [9:0]  io_col,
  input  [7:0]  io_in_0,
  input  [7:0]  io_in_1,
  input  [7:0]  io_in_2,
  input  [7:0]  io_in_3,
  input  [7:0]  io_in_4,
  input  [7:0]  io_in_5,
  input  [7:0]  io_in_6,
  input  [7:0]  io_in_7,
  output [31:0] io_ifm_o_data_0,
  output [31:0] io_ifm_o_data_1,
  output [31:0] io_ifm_o_data_2,
  output [31:0] io_ifm_o_data_3,
  output [31:0] io_ifm_o_data_4,
  output [31:0] io_ifm_o_data_5,
  output [31:0] io_ifm_o_data_6,
  output [31:0] io_ifm_o_data_7,
  input         io_pad_top,
  input         io_pad_bottom,
  input         io_pad_left_and_right,
  input  [4:0]  io_zero_pad_valid_s2,
  input         io_zero_pad_valid_s1,
  input  [7:0]  io_zero_point_in
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
`endif // RANDOMIZE_REG_INIT
  wire  TPRAM_WRAP_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_1_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_1_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_1_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_1_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_2_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_2_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_2_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_2_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_3_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_3_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_3_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_3_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_4_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_4_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_4_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_4_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_5_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_5_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_5_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_5_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_6_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_6_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_6_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_6_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_7_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_7_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_7_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_7_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_8_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_8_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_8_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_8_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_8_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_8_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_8_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_9_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_9_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_9_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_9_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_9_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_9_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_9_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_10_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_10_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_10_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_10_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_10_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_10_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_10_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_11_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_11_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_11_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_11_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_11_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_11_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_11_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_12_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_12_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_12_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_12_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_12_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_12_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_12_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_13_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_13_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_13_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_13_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_13_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_13_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_13_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_14_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_14_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_14_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_14_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_14_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_14_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_14_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_15_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_15_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_15_io_ren; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_15_io_waddr; // @[utils.scala 237:100]
  wire [10:0] TPRAM_WRAP_15_io_raddr; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_15_io_wdata; // @[utils.scala 237:100]
  wire [15:0] TPRAM_WRAP_15_io_rdata; // @[utils.scala 237:100]
  reg  in_temp_sel; // @[IfmBuffer.scala 42:30]
  wire  _in_temp_sel_T = ~in_temp_sel; // @[IfmBuffer.scala 43:67]
  reg [7:0] in_temp_0; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_1; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_2; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_3; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_4; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_5; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_6; // @[IfmBuffer.scala 44:39]
  reg [7:0] in_temp_7; // @[IfmBuffer.scala 44:39]
  wire [15:0] _write_data_0_T = {io_in_0,io_in_0}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_0_T_1 = {io_in_0,in_temp_0}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_1_T = {io_in_1,io_in_1}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_1_T_1 = {io_in_1,in_temp_1}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_2_T = {io_in_2,io_in_2}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_2_T_1 = {io_in_2,in_temp_2}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_3_T = {io_in_3,io_in_3}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_3_T_1 = {io_in_3,in_temp_3}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_4_T = {io_in_4,io_in_4}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_4_T_1 = {io_in_4,in_temp_4}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_5_T = {io_in_5,io_in_5}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_5_T_1 = {io_in_5,in_temp_5}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_6_T = {io_in_6,io_in_6}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_6_T_1 = {io_in_6,in_temp_6}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_7_T = {io_in_7,io_in_7}; // @[Cat.scala 33:92]
  wire [15:0] _write_data_7_T_1 = {io_in_7,in_temp_7}; // @[Cat.scala 33:92]
  reg  row_is_singal_or_double; // @[IfmBuffer.scala 52:40]
  reg [9:0] col_cnt; // @[IfmBuffer.scala 55:24]
  wire [9:0] _col_cnt_T_1 = io_col - 10'h1; // @[IfmBuffer.scala 56:77]
  wire  _col_cnt_T_2 = col_cnt == _col_cnt_T_1; // @[IfmBuffer.scala 56:67]
  wire [9:0] _col_cnt_T_4 = col_cnt + 10'h1; // @[IfmBuffer.scala 56:94]
  wire  _row_is_singal_or_double_T_3 = ~row_is_singal_or_double; // @[IfmBuffer.scala 57:89]
  reg [10:0] bram_write_addr_singal; // @[IfmBuffer.scala 62:40]
  reg [10:0] bram_write_addr_double; // @[IfmBuffer.scala 63:41]
  wire [10:0] _bram_write_addr_singal_T_2 = bram_write_addr_singal + 11'h1; // @[IfmBuffer.scala 64:107]
  wire [11:0] _GEN_2 = {{1'd0}, _bram_write_addr_singal_T_2}; // @[IfmBuffer.scala 64:111]
  wire [11:0] _bram_write_addr_singal_T_3 = _GEN_2 << io_upsample_enable; // @[IfmBuffer.scala 64:111]
  wire [11:0] _bram_write_addr_singal_T_4 = io_bram_en_write & _row_is_singal_or_double_T_3 ?
    _bram_write_addr_singal_T_3 : {{1'd0}, bram_write_addr_singal}; // @[IfmBuffer.scala 64:53]
  wire [11:0] _bram_write_addr_singal_T_5 = io_recv_done ? 12'h0 : _bram_write_addr_singal_T_4; // @[IfmBuffer.scala 64:32]
  wire [10:0] _bram_write_addr_double_T_2 = bram_write_addr_double + 11'h1; // @[IfmBuffer.scala 65:107]
  wire [11:0] _GEN_3 = {{1'd0}, _bram_write_addr_double_T_2}; // @[IfmBuffer.scala 65:111]
  wire [11:0] _bram_write_addr_double_T_3 = _GEN_3 << io_upsample_enable; // @[IfmBuffer.scala 65:111]
  wire [11:0] _bram_write_addr_double_T_4 = io_bram_en_write & row_is_singal_or_double ? _bram_write_addr_double_T_3 :
    {{1'd0}, bram_write_addr_double}; // @[IfmBuffer.scala 65:53]
  wire [11:0] _bram_write_addr_double_T_5 = io_recv_done ? 12'h0 : _bram_write_addr_double_T_4; // @[IfmBuffer.scala 65:32]
  wire  read_singal_row_s1 = ~io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 67:87]
  wire [9:0] bram_read_addr_singal = io_ifmbuf_bram_addr_read_s1[9:0]; // @[IfmBuffer.scala 69:58]
  wire  _bram_read_addr_s1_singal_extend_T = ~io_buf_sel; // @[IfmBuffer.scala 74:46]
  wire [10:0] bram_read_addr_s1_singal_extend = {_bram_read_addr_s1_singal_extend_T,bram_read_addr_singal}; // @[Cat.scala 33:92]
  wire [10:0] bram_read_addr_s2_singal_extend = {_bram_read_addr_s1_singal_extend_T,io_ifmbuf_bram_addr_read_s2_singal}; // @[Cat.scala 33:92]
  wire [10:0] bram_read_addr_s2_double_extend = {_bram_read_addr_s1_singal_extend_T,io_ifmbuf_bram_addr_read_s2_double}; // @[Cat.scala 33:92]
  wire [15:0] temp_single_0 = TPRAM_WRAP_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_0_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_0 = TPRAM_WRAP_8_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_0_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_1 = TPRAM_WRAP_1_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_1_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_1 = TPRAM_WRAP_9_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_1_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_2 = TPRAM_WRAP_2_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_2_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_2 = TPRAM_WRAP_10_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_2_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_3 = TPRAM_WRAP_3_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_3_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_3 = TPRAM_WRAP_11_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_3_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_4 = TPRAM_WRAP_4_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_4_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_4 = TPRAM_WRAP_12_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_4_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_5 = TPRAM_WRAP_5_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_5_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_5 = TPRAM_WRAP_13_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_5_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_6 = TPRAM_WRAP_6_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_6_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_6 = TPRAM_WRAP_14_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_6_REG; // @[IfmBuffer.scala 85:40]
  wire [15:0] temp_single_7 = TPRAM_WRAP_7_io_rdata; // @[IfmBuffer.scala 79:27 97:24]
  reg [7:0] temp_single_regnext_7_REG; // @[IfmBuffer.scala 84:40]
  wire [15:0] temp_double_7 = TPRAM_WRAP_15_io_rdata; // @[IfmBuffer.scala 104:24 80:27]
  reg [7:0] temp_double_regnext_7_REG; // @[IfmBuffer.scala 85:40]
  wire  _T_1 = io_bram_en_write & (in_temp_sel | io_upsample_enable); // @[IfmBuffer.scala 92:47]
  wire  _T_3 = ~io_s_mod; // @[IfmBuffer.scala 93:43]
  wire  zero_s2_pad_left = io_zero_pad_valid_s2[4]; // @[IfmBuffer.scala 110:48]
  wire  zero_s2_pad_right = io_zero_pad_valid_s2[3]; // @[IfmBuffer.scala 111:49]
  wire  zero_s2_pad_top = io_zero_pad_valid_s2[2]; // @[IfmBuffer.scala 112:47]
  wire  zero_s2_pad_only_bottom = io_zero_pad_valid_s2[1]; // @[IfmBuffer.scala 113:55]
  wire  zero_s2_pad_bottom_include_top = io_zero_pad_valid_s2[0]; // @[IfmBuffer.scala 114:62]
  wire  pad_require = io_pad_top | io_pad_bottom | io_pad_left_and_right; // @[IfmBuffer.scala 129:48]
  wire [7:0] out_s1_singal_0 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_0[15:8] : temp_single_0[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_0 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_0[15:8] : temp_double_0[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_0_T = read_singal_row_s1 ? out_s1_singal_0 : out_s1_double_0; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_0 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_0_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_0_T_1 = {temp_single_0[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_0_T_2 = {io_zero_point_in,temp_single_regnext_0_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_0_T_4 = {temp_single_0[7:0],temp_single_regnext_0_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_0_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_0_T_2 :
    _out_s2_pad_left_and_right_signal_0_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_0 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_0_T_1 :
    _out_s2_pad_left_and_right_signal_0_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_0_T_1 = {temp_double_0[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_0_T_2 = {io_zero_point_in,temp_double_regnext_0_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_0_T_4 = {temp_double_0[7:0],temp_double_regnext_0_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_0_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_0_T_2 :
    _out_s2_pad_left_and_right_double_0_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_0 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_0_T_1 :
    _out_s2_pad_left_and_right_double_0_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_0_T_1 = {out_s2_pad_left_and_right_signal_0,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_0_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_0}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_0_T_4 = {out_s2_pad_left_and_right_signal_0,
    out_s2_pad_left_and_right_double_0}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_0_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_0_T_3 : _out_s2_pad_top_however_bottom_0_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_0 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_0_T_1 :
    _out_s2_pad_top_however_bottom_0_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_0_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_0}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_0_T_2 = {out_s2_pad_left_and_right_double_0,out_s2_pad_left_and_right_signal_0}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_0 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_0_T_1 :
    _out_s2_pad_only_bottom_0_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_0_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_0 : _out_s2_pad_only_bottom_0_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_0 = io_pad_top ? out_s2_pad_top_however_bottom_0 : _out_s2_pad_0_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_0_T = {temp_double_0,temp_single_0}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_0 = pad_require ? out_s2_pad_0 : _out_s2_0_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_0_T = {24'h0,out_s1_0}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_1 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_1[15:8] : temp_single_1[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_1 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_1[15:8] : temp_double_1[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_1_T = read_singal_row_s1 ? out_s1_singal_1 : out_s1_double_1; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_1 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_1_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_1_T_1 = {temp_single_1[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_1_T_2 = {io_zero_point_in,temp_single_regnext_1_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_1_T_4 = {temp_single_1[7:0],temp_single_regnext_1_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_1_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_1_T_2 :
    _out_s2_pad_left_and_right_signal_1_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_1 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_1_T_1 :
    _out_s2_pad_left_and_right_signal_1_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_1_T_1 = {temp_double_1[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_1_T_2 = {io_zero_point_in,temp_double_regnext_1_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_1_T_4 = {temp_double_1[7:0],temp_double_regnext_1_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_1_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_1_T_2 :
    _out_s2_pad_left_and_right_double_1_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_1 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_1_T_1 :
    _out_s2_pad_left_and_right_double_1_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_1_T_1 = {out_s2_pad_left_and_right_signal_1,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_1_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_1}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_1_T_4 = {out_s2_pad_left_and_right_signal_1,
    out_s2_pad_left_and_right_double_1}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_1_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_1_T_3 : _out_s2_pad_top_however_bottom_1_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_1 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_1_T_1 :
    _out_s2_pad_top_however_bottom_1_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_1_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_1}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_1_T_2 = {out_s2_pad_left_and_right_double_1,out_s2_pad_left_and_right_signal_1}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_1 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_1_T_1 :
    _out_s2_pad_only_bottom_1_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_1_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_1 : _out_s2_pad_only_bottom_1_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_1 = io_pad_top ? out_s2_pad_top_however_bottom_1 : _out_s2_pad_1_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_1_T = {temp_double_1,temp_single_1}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_1 = pad_require ? out_s2_pad_1 : _out_s2_1_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_1_T = {24'h0,out_s1_1}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_2 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_2[15:8] : temp_single_2[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_2 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_2[15:8] : temp_double_2[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_2_T = read_singal_row_s1 ? out_s1_singal_2 : out_s1_double_2; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_2 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_2_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_2_T_1 = {temp_single_2[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_2_T_2 = {io_zero_point_in,temp_single_regnext_2_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_2_T_4 = {temp_single_2[7:0],temp_single_regnext_2_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_2_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_2_T_2 :
    _out_s2_pad_left_and_right_signal_2_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_2 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_2_T_1 :
    _out_s2_pad_left_and_right_signal_2_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_2_T_1 = {temp_double_2[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_2_T_2 = {io_zero_point_in,temp_double_regnext_2_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_2_T_4 = {temp_double_2[7:0],temp_double_regnext_2_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_2_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_2_T_2 :
    _out_s2_pad_left_and_right_double_2_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_2 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_2_T_1 :
    _out_s2_pad_left_and_right_double_2_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_2_T_1 = {out_s2_pad_left_and_right_signal_2,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_2_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_2}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_2_T_4 = {out_s2_pad_left_and_right_signal_2,
    out_s2_pad_left_and_right_double_2}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_2_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_2_T_3 : _out_s2_pad_top_however_bottom_2_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_2 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_2_T_1 :
    _out_s2_pad_top_however_bottom_2_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_2_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_2}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_2_T_2 = {out_s2_pad_left_and_right_double_2,out_s2_pad_left_and_right_signal_2}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_2 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_2_T_1 :
    _out_s2_pad_only_bottom_2_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_2_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_2 : _out_s2_pad_only_bottom_2_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_2 = io_pad_top ? out_s2_pad_top_however_bottom_2 : _out_s2_pad_2_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_2_T = {temp_double_2,temp_single_2}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_2 = pad_require ? out_s2_pad_2 : _out_s2_2_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_2_T = {24'h0,out_s1_2}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_3 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_3[15:8] : temp_single_3[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_3 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_3[15:8] : temp_double_3[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_3_T = read_singal_row_s1 ? out_s1_singal_3 : out_s1_double_3; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_3 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_3_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_3_T_1 = {temp_single_3[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_3_T_2 = {io_zero_point_in,temp_single_regnext_3_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_3_T_4 = {temp_single_3[7:0],temp_single_regnext_3_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_3_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_3_T_2 :
    _out_s2_pad_left_and_right_signal_3_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_3 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_3_T_1 :
    _out_s2_pad_left_and_right_signal_3_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_3_T_1 = {temp_double_3[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_3_T_2 = {io_zero_point_in,temp_double_regnext_3_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_3_T_4 = {temp_double_3[7:0],temp_double_regnext_3_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_3_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_3_T_2 :
    _out_s2_pad_left_and_right_double_3_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_3 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_3_T_1 :
    _out_s2_pad_left_and_right_double_3_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_3_T_1 = {out_s2_pad_left_and_right_signal_3,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_3_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_3}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_3_T_4 = {out_s2_pad_left_and_right_signal_3,
    out_s2_pad_left_and_right_double_3}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_3_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_3_T_3 : _out_s2_pad_top_however_bottom_3_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_3 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_3_T_1 :
    _out_s2_pad_top_however_bottom_3_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_3_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_3}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_3_T_2 = {out_s2_pad_left_and_right_double_3,out_s2_pad_left_and_right_signal_3}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_3 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_3_T_1 :
    _out_s2_pad_only_bottom_3_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_3_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_3 : _out_s2_pad_only_bottom_3_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_3 = io_pad_top ? out_s2_pad_top_however_bottom_3 : _out_s2_pad_3_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_3_T = {temp_double_3,temp_single_3}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_3 = pad_require ? out_s2_pad_3 : _out_s2_3_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_3_T = {24'h0,out_s1_3}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_4 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_4[15:8] : temp_single_4[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_4 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_4[15:8] : temp_double_4[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_4_T = read_singal_row_s1 ? out_s1_singal_4 : out_s1_double_4; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_4 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_4_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_4_T_1 = {temp_single_4[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_4_T_2 = {io_zero_point_in,temp_single_regnext_4_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_4_T_4 = {temp_single_4[7:0],temp_single_regnext_4_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_4_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_4_T_2 :
    _out_s2_pad_left_and_right_signal_4_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_4 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_4_T_1 :
    _out_s2_pad_left_and_right_signal_4_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_4_T_1 = {temp_double_4[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_4_T_2 = {io_zero_point_in,temp_double_regnext_4_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_4_T_4 = {temp_double_4[7:0],temp_double_regnext_4_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_4_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_4_T_2 :
    _out_s2_pad_left_and_right_double_4_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_4 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_4_T_1 :
    _out_s2_pad_left_and_right_double_4_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_4_T_1 = {out_s2_pad_left_and_right_signal_4,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_4_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_4}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_4_T_4 = {out_s2_pad_left_and_right_signal_4,
    out_s2_pad_left_and_right_double_4}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_4_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_4_T_3 : _out_s2_pad_top_however_bottom_4_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_4 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_4_T_1 :
    _out_s2_pad_top_however_bottom_4_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_4_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_4}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_4_T_2 = {out_s2_pad_left_and_right_double_4,out_s2_pad_left_and_right_signal_4}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_4 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_4_T_1 :
    _out_s2_pad_only_bottom_4_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_4_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_4 : _out_s2_pad_only_bottom_4_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_4 = io_pad_top ? out_s2_pad_top_however_bottom_4 : _out_s2_pad_4_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_4_T = {temp_double_4,temp_single_4}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_4 = pad_require ? out_s2_pad_4 : _out_s2_4_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_4_T = {24'h0,out_s1_4}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_5 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_5[15:8] : temp_single_5[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_5 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_5[15:8] : temp_double_5[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_5_T = read_singal_row_s1 ? out_s1_singal_5 : out_s1_double_5; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_5 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_5_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_5_T_1 = {temp_single_5[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_5_T_2 = {io_zero_point_in,temp_single_regnext_5_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_5_T_4 = {temp_single_5[7:0],temp_single_regnext_5_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_5_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_5_T_2 :
    _out_s2_pad_left_and_right_signal_5_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_5 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_5_T_1 :
    _out_s2_pad_left_and_right_signal_5_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_5_T_1 = {temp_double_5[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_5_T_2 = {io_zero_point_in,temp_double_regnext_5_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_5_T_4 = {temp_double_5[7:0],temp_double_regnext_5_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_5_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_5_T_2 :
    _out_s2_pad_left_and_right_double_5_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_5 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_5_T_1 :
    _out_s2_pad_left_and_right_double_5_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_5_T_1 = {out_s2_pad_left_and_right_signal_5,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_5_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_5}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_5_T_4 = {out_s2_pad_left_and_right_signal_5,
    out_s2_pad_left_and_right_double_5}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_5_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_5_T_3 : _out_s2_pad_top_however_bottom_5_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_5 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_5_T_1 :
    _out_s2_pad_top_however_bottom_5_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_5_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_5}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_5_T_2 = {out_s2_pad_left_and_right_double_5,out_s2_pad_left_and_right_signal_5}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_5 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_5_T_1 :
    _out_s2_pad_only_bottom_5_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_5_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_5 : _out_s2_pad_only_bottom_5_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_5 = io_pad_top ? out_s2_pad_top_however_bottom_5 : _out_s2_pad_5_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_5_T = {temp_double_5,temp_single_5}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_5 = pad_require ? out_s2_pad_5 : _out_s2_5_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_5_T = {24'h0,out_s1_5}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_6 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_6[15:8] : temp_single_6[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_6 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_6[15:8] : temp_double_6[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_6_T = read_singal_row_s1 ? out_s1_singal_6 : out_s1_double_6; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_6 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_6_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_6_T_1 = {temp_single_6[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_6_T_2 = {io_zero_point_in,temp_single_regnext_6_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_6_T_4 = {temp_single_6[7:0],temp_single_regnext_6_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_6_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_6_T_2 :
    _out_s2_pad_left_and_right_signal_6_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_6 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_6_T_1 :
    _out_s2_pad_left_and_right_signal_6_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_6_T_1 = {temp_double_6[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_6_T_2 = {io_zero_point_in,temp_double_regnext_6_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_6_T_4 = {temp_double_6[7:0],temp_double_regnext_6_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_6_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_6_T_2 :
    _out_s2_pad_left_and_right_double_6_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_6 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_6_T_1 :
    _out_s2_pad_left_and_right_double_6_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_6_T_1 = {out_s2_pad_left_and_right_signal_6,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_6_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_6}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_6_T_4 = {out_s2_pad_left_and_right_signal_6,
    out_s2_pad_left_and_right_double_6}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_6_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_6_T_3 : _out_s2_pad_top_however_bottom_6_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_6 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_6_T_1 :
    _out_s2_pad_top_however_bottom_6_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_6_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_6}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_6_T_2 = {out_s2_pad_left_and_right_double_6,out_s2_pad_left_and_right_signal_6}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_6 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_6_T_1 :
    _out_s2_pad_only_bottom_6_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_6_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_6 : _out_s2_pad_only_bottom_6_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_6 = io_pad_top ? out_s2_pad_top_however_bottom_6 : _out_s2_pad_6_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_6_T = {temp_double_6,temp_single_6}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_6 = pad_require ? out_s2_pad_6 : _out_s2_6_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_6_T = {24'h0,out_s1_6}; // @[Cat.scala 33:92]
  wire [7:0] out_s1_singal_7 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_single_7[15:8] : temp_single_7[7:0]; // @[IfmBuffer.scala 132:30]
  wire [7:0] out_s1_double_7 = io_ifmbuf_bram_addr_read_sel_s1 ? temp_double_7[15:8] : temp_double_7[7:0]; // @[IfmBuffer.scala 133:30]
  wire [7:0] _out_s1_7_T = read_singal_row_s1 ? out_s1_singal_7 : out_s1_double_7; // @[IfmBuffer.scala 135:58]
  wire [7:0] out_s1_7 = io_zero_pad_valid_s1 ? io_zero_point_in : _out_s1_7_T; // @[IfmBuffer.scala 135:23]
  wire [15:0] _out_s2_pad_left_and_right_signal_7_T_1 = {temp_single_7[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_7_T_2 = {io_zero_point_in,temp_single_regnext_7_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_7_T_4 = {temp_single_7[7:0],temp_single_regnext_7_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_signal_7_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_signal_7_T_2 :
    _out_s2_pad_left_and_right_signal_7_T_4; // @[IfmBuffer.scala 137:115]
  wire [15:0] out_s2_pad_left_and_right_signal_7 = zero_s2_pad_left ? _out_s2_pad_left_and_right_signal_7_T_1 :
    _out_s2_pad_left_and_right_signal_7_T_5; // @[IfmBuffer.scala 137:49]
  wire [15:0] _out_s2_pad_left_and_right_double_7_T_1 = {temp_double_7[7:0],io_zero_point_in}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_7_T_2 = {io_zero_point_in,temp_double_regnext_7_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_7_T_4 = {temp_double_7[7:0],temp_double_regnext_7_REG}; // @[Cat.scala 33:92]
  wire [15:0] _out_s2_pad_left_and_right_double_7_T_5 = zero_s2_pad_right ? _out_s2_pad_left_and_right_double_7_T_2 :
    _out_s2_pad_left_and_right_double_7_T_4; // @[IfmBuffer.scala 138:115]
  wire [15:0] out_s2_pad_left_and_right_double_7 = zero_s2_pad_left ? _out_s2_pad_left_and_right_double_7_T_1 :
    _out_s2_pad_left_and_right_double_7_T_5; // @[IfmBuffer.scala 138:49]
  wire [31:0] _out_s2_pad_top_however_bottom_7_T_1 = {out_s2_pad_left_and_right_signal_7,io_zero_point_in,
    io_zero_point_in}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_7_T_3 = {io_zero_point_in,io_zero_point_in,
    out_s2_pad_left_and_right_double_7}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_7_T_4 = {out_s2_pad_left_and_right_signal_7,
    out_s2_pad_left_and_right_double_7}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_top_however_bottom_7_T_5 = zero_s2_pad_bottom_include_top ?
    _out_s2_pad_top_however_bottom_7_T_3 : _out_s2_pad_top_however_bottom_7_T_4; // @[IfmBuffer.scala 139:125]
  wire [31:0] out_s2_pad_top_however_bottom_7 = zero_s2_pad_top ? _out_s2_pad_top_however_bottom_7_T_1 :
    _out_s2_pad_top_however_bottom_7_T_5; // @[IfmBuffer.scala 139:46]
  wire [31:0] _out_s2_pad_only_bottom_7_T_1 = {io_zero_point_in,io_zero_point_in,out_s2_pad_left_and_right_signal_7}; // @[Cat.scala 33:92]
  wire [31:0] _out_s2_pad_only_bottom_7_T_2 = {out_s2_pad_left_and_right_double_7,out_s2_pad_left_and_right_signal_7}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_pad_only_bottom_7 = zero_s2_pad_only_bottom ? _out_s2_pad_only_bottom_7_T_1 :
    _out_s2_pad_only_bottom_7_T_2; // @[IfmBuffer.scala 140:39]
  wire [31:0] _out_s2_pad_7_T_1 = io_pad_bottom ? out_s2_pad_only_bottom_7 : _out_s2_pad_only_bottom_7_T_2; // @[IfmBuffer.scala 141:75]
  wire [31:0] out_s2_pad_7 = io_pad_top ? out_s2_pad_top_however_bottom_7 : _out_s2_pad_7_T_1; // @[IfmBuffer.scala 141:27]
  wire [31:0] _out_s2_7_T = {temp_double_7,temp_single_7}; // @[Cat.scala 33:92]
  wire [31:0] out_s2_7 = pad_require ? out_s2_pad_7 : _out_s2_7_T; // @[IfmBuffer.scala 142:23]
  wire [31:0] _io_ifm_o_data_7_T = {24'h0,out_s1_7}; // @[Cat.scala 33:92]
  wire [11:0] _GEN_0 = reset ? 12'h0 : _bram_write_addr_singal_T_5; // @[IfmBuffer.scala 62:{40,40} 64:27]
  wire [11:0] _GEN_1 = reset ? 12'h0 : _bram_write_addr_double_T_5; // @[IfmBuffer.scala 63:{41,41} 65:27]
  TPRAM_WRAP TPRAM_WRAP ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_clock),
    .io_wen(TPRAM_WRAP_io_wen),
    .io_ren(TPRAM_WRAP_io_ren),
    .io_waddr(TPRAM_WRAP_io_waddr),
    .io_raddr(TPRAM_WRAP_io_raddr),
    .io_wdata(TPRAM_WRAP_io_wdata),
    .io_rdata(TPRAM_WRAP_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_1 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_1_clock),
    .io_wen(TPRAM_WRAP_1_io_wen),
    .io_ren(TPRAM_WRAP_1_io_ren),
    .io_waddr(TPRAM_WRAP_1_io_waddr),
    .io_raddr(TPRAM_WRAP_1_io_raddr),
    .io_wdata(TPRAM_WRAP_1_io_wdata),
    .io_rdata(TPRAM_WRAP_1_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_2 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_2_clock),
    .io_wen(TPRAM_WRAP_2_io_wen),
    .io_ren(TPRAM_WRAP_2_io_ren),
    .io_waddr(TPRAM_WRAP_2_io_waddr),
    .io_raddr(TPRAM_WRAP_2_io_raddr),
    .io_wdata(TPRAM_WRAP_2_io_wdata),
    .io_rdata(TPRAM_WRAP_2_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_3 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_3_clock),
    .io_wen(TPRAM_WRAP_3_io_wen),
    .io_ren(TPRAM_WRAP_3_io_ren),
    .io_waddr(TPRAM_WRAP_3_io_waddr),
    .io_raddr(TPRAM_WRAP_3_io_raddr),
    .io_wdata(TPRAM_WRAP_3_io_wdata),
    .io_rdata(TPRAM_WRAP_3_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_4 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_4_clock),
    .io_wen(TPRAM_WRAP_4_io_wen),
    .io_ren(TPRAM_WRAP_4_io_ren),
    .io_waddr(TPRAM_WRAP_4_io_waddr),
    .io_raddr(TPRAM_WRAP_4_io_raddr),
    .io_wdata(TPRAM_WRAP_4_io_wdata),
    .io_rdata(TPRAM_WRAP_4_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_5 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_5_clock),
    .io_wen(TPRAM_WRAP_5_io_wen),
    .io_ren(TPRAM_WRAP_5_io_ren),
    .io_waddr(TPRAM_WRAP_5_io_waddr),
    .io_raddr(TPRAM_WRAP_5_io_raddr),
    .io_wdata(TPRAM_WRAP_5_io_wdata),
    .io_rdata(TPRAM_WRAP_5_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_6 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_6_clock),
    .io_wen(TPRAM_WRAP_6_io_wen),
    .io_ren(TPRAM_WRAP_6_io_ren),
    .io_waddr(TPRAM_WRAP_6_io_waddr),
    .io_raddr(TPRAM_WRAP_6_io_raddr),
    .io_wdata(TPRAM_WRAP_6_io_wdata),
    .io_rdata(TPRAM_WRAP_6_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_7 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_7_clock),
    .io_wen(TPRAM_WRAP_7_io_wen),
    .io_ren(TPRAM_WRAP_7_io_ren),
    .io_waddr(TPRAM_WRAP_7_io_waddr),
    .io_raddr(TPRAM_WRAP_7_io_raddr),
    .io_wdata(TPRAM_WRAP_7_io_wdata),
    .io_rdata(TPRAM_WRAP_7_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_8 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_8_clock),
    .io_wen(TPRAM_WRAP_8_io_wen),
    .io_ren(TPRAM_WRAP_8_io_ren),
    .io_waddr(TPRAM_WRAP_8_io_waddr),
    .io_raddr(TPRAM_WRAP_8_io_raddr),
    .io_wdata(TPRAM_WRAP_8_io_wdata),
    .io_rdata(TPRAM_WRAP_8_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_9 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_9_clock),
    .io_wen(TPRAM_WRAP_9_io_wen),
    .io_ren(TPRAM_WRAP_9_io_ren),
    .io_waddr(TPRAM_WRAP_9_io_waddr),
    .io_raddr(TPRAM_WRAP_9_io_raddr),
    .io_wdata(TPRAM_WRAP_9_io_wdata),
    .io_rdata(TPRAM_WRAP_9_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_10 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_10_clock),
    .io_wen(TPRAM_WRAP_10_io_wen),
    .io_ren(TPRAM_WRAP_10_io_ren),
    .io_waddr(TPRAM_WRAP_10_io_waddr),
    .io_raddr(TPRAM_WRAP_10_io_raddr),
    .io_wdata(TPRAM_WRAP_10_io_wdata),
    .io_rdata(TPRAM_WRAP_10_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_11 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_11_clock),
    .io_wen(TPRAM_WRAP_11_io_wen),
    .io_ren(TPRAM_WRAP_11_io_ren),
    .io_waddr(TPRAM_WRAP_11_io_waddr),
    .io_raddr(TPRAM_WRAP_11_io_raddr),
    .io_wdata(TPRAM_WRAP_11_io_wdata),
    .io_rdata(TPRAM_WRAP_11_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_12 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_12_clock),
    .io_wen(TPRAM_WRAP_12_io_wen),
    .io_ren(TPRAM_WRAP_12_io_ren),
    .io_waddr(TPRAM_WRAP_12_io_waddr),
    .io_raddr(TPRAM_WRAP_12_io_raddr),
    .io_wdata(TPRAM_WRAP_12_io_wdata),
    .io_rdata(TPRAM_WRAP_12_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_13 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_13_clock),
    .io_wen(TPRAM_WRAP_13_io_wen),
    .io_ren(TPRAM_WRAP_13_io_ren),
    .io_waddr(TPRAM_WRAP_13_io_waddr),
    .io_raddr(TPRAM_WRAP_13_io_raddr),
    .io_wdata(TPRAM_WRAP_13_io_wdata),
    .io_rdata(TPRAM_WRAP_13_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_14 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_14_clock),
    .io_wen(TPRAM_WRAP_14_io_wen),
    .io_ren(TPRAM_WRAP_14_io_ren),
    .io_waddr(TPRAM_WRAP_14_io_waddr),
    .io_raddr(TPRAM_WRAP_14_io_raddr),
    .io_wdata(TPRAM_WRAP_14_io_wdata),
    .io_rdata(TPRAM_WRAP_14_io_rdata)
  );
  TPRAM_WRAP TPRAM_WRAP_15 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_15_clock),
    .io_wen(TPRAM_WRAP_15_io_wen),
    .io_ren(TPRAM_WRAP_15_io_ren),
    .io_waddr(TPRAM_WRAP_15_io_waddr),
    .io_raddr(TPRAM_WRAP_15_io_raddr),
    .io_wdata(TPRAM_WRAP_15_io_wdata),
    .io_rdata(TPRAM_WRAP_15_io_rdata)
  );
  assign io_ifm_o_data_0 = io_s_mod ? out_s2_0 : _io_ifm_o_data_0_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_1 = io_s_mod ? out_s2_1 : _io_ifm_o_data_1_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_2 = io_s_mod ? out_s2_2 : _io_ifm_o_data_2_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_3 = io_s_mod ? out_s2_3 : _io_ifm_o_data_3_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_4 = io_s_mod ? out_s2_4 : _io_ifm_o_data_4_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_5 = io_s_mod ? out_s2_5 : _io_ifm_o_data_5_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_6 = io_s_mod ? out_s2_6 : _io_ifm_o_data_6_T; // @[IfmBuffer.scala 144:30]
  assign io_ifm_o_data_7 = io_s_mod ? out_s2_7 : _io_ifm_o_data_7_T; // @[IfmBuffer.scala 144:30]
  assign TPRAM_WRAP_clock = clock;
  assign TPRAM_WRAP_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_io_wdata = io_upsample_enable ? _write_data_0_T : _write_data_0_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_1_clock = clock;
  assign TPRAM_WRAP_1_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_1_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_1_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_1_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_1_io_wdata = io_upsample_enable ? _write_data_1_T : _write_data_1_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_2_clock = clock;
  assign TPRAM_WRAP_2_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_2_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_2_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_2_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_2_io_wdata = io_upsample_enable ? _write_data_2_T : _write_data_2_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_3_clock = clock;
  assign TPRAM_WRAP_3_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_3_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_3_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_3_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_3_io_wdata = io_upsample_enable ? _write_data_3_T : _write_data_3_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_4_clock = clock;
  assign TPRAM_WRAP_4_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_4_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_4_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_4_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_4_io_wdata = io_upsample_enable ? _write_data_4_T : _write_data_4_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_5_clock = clock;
  assign TPRAM_WRAP_5_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_5_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_5_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_5_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_5_io_wdata = io_upsample_enable ? _write_data_5_T : _write_data_5_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_6_clock = clock;
  assign TPRAM_WRAP_6_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_6_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_6_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_6_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_6_io_wdata = io_upsample_enable ? _write_data_6_T : _write_data_6_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_7_clock = clock;
  assign TPRAM_WRAP_7_io_wen = io_bram_en_write & (in_temp_sel | io_upsample_enable) & _row_is_singal_or_double_T_3; // @[IfmBuffer.scala 92:83]
  assign TPRAM_WRAP_7_io_ren = io_s_mod | ~io_s_mod & read_singal_row_s1; // @[IfmBuffer.scala 93:39]
  assign TPRAM_WRAP_7_io_waddr = {io_buf_sel,bram_write_addr_singal[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_7_io_raddr = io_s_mod ? bram_read_addr_s2_singal_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 95:35]
  assign TPRAM_WRAP_7_io_wdata = io_upsample_enable ? _write_data_7_T : _write_data_7_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_8_clock = clock;
  assign TPRAM_WRAP_8_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_8_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_8_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_8_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_8_io_wdata = io_upsample_enable ? _write_data_0_T : _write_data_0_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_9_clock = clock;
  assign TPRAM_WRAP_9_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_9_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_9_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_9_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_9_io_wdata = io_upsample_enable ? _write_data_1_T : _write_data_1_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_10_clock = clock;
  assign TPRAM_WRAP_10_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_10_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_10_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_10_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_10_io_wdata = io_upsample_enable ? _write_data_2_T : _write_data_2_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_11_clock = clock;
  assign TPRAM_WRAP_11_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_11_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_11_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_11_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_11_io_wdata = io_upsample_enable ? _write_data_3_T : _write_data_3_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_12_clock = clock;
  assign TPRAM_WRAP_12_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_12_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_12_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_12_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_12_io_wdata = io_upsample_enable ? _write_data_4_T : _write_data_4_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_13_clock = clock;
  assign TPRAM_WRAP_13_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_13_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_13_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_13_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_13_io_wdata = io_upsample_enable ? _write_data_5_T : _write_data_5_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_14_clock = clock;
  assign TPRAM_WRAP_14_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_14_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_14_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_14_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_14_io_wdata = io_upsample_enable ? _write_data_6_T : _write_data_6_T_1; // @[IfmBuffer.scala 48:29]
  assign TPRAM_WRAP_15_clock = clock;
  assign TPRAM_WRAP_15_io_wen = _T_1 & row_is_singal_or_double; // @[IfmBuffer.scala 99:83]
  assign TPRAM_WRAP_15_io_ren = io_s_mod | _T_3 & io_ifmbuf_bram_addr_read_s1[10]; // @[IfmBuffer.scala 100:39]
  assign TPRAM_WRAP_15_io_waddr = {io_buf_sel,bram_write_addr_double[10:1]}; // @[Cat.scala 33:92]
  assign TPRAM_WRAP_15_io_raddr = io_s_mod ? bram_read_addr_s2_double_extend : bram_read_addr_s1_singal_extend; // @[IfmBuffer.scala 102:35]
  assign TPRAM_WRAP_15_io_wdata = io_upsample_enable ? _write_data_7_T : _write_data_7_T_1; // @[IfmBuffer.scala 48:29]
  always @(posedge clock) begin
    if (reset) begin // @[IfmBuffer.scala 42:30]
      in_temp_sel <= 1'h0; // @[IfmBuffer.scala 42:30]
    end else if (io_recv_done) begin // @[IfmBuffer.scala 43:23]
      in_temp_sel <= 1'h0;
    end else if (io_bram_en_write) begin // @[IfmBuffer.scala 43:48]
      in_temp_sel <= ~in_temp_sel;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_0 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_0 <= io_in_0;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_1 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_1 <= io_in_1;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_2 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_2 <= io_in_2;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_3 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_3 <= io_in_3;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_4 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_4 <= io_in_4;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_5 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_5 <= io_in_5;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_6 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_6 <= io_in_6;
    end
    if (reset) begin // @[IfmBuffer.scala 44:39]
      in_temp_7 <= 8'h0; // @[IfmBuffer.scala 44:39]
    end else if (_in_temp_sel_T) begin // @[IfmBuffer.scala 47:24]
      in_temp_7 <= io_in_7;
    end
    if (reset) begin // @[IfmBuffer.scala 52:40]
      row_is_singal_or_double <= 1'h0; // @[IfmBuffer.scala 52:40]
    end else if (io_recv_done) begin // @[IfmBuffer.scala 57:35]
      row_is_singal_or_double <= 1'h0;
    end else if (_col_cnt_T_2) begin // @[IfmBuffer.scala 57:60]
      row_is_singal_or_double <= ~row_is_singal_or_double;
    end
    if (reset) begin // @[IfmBuffer.scala 55:24]
      col_cnt <= 10'h0; // @[IfmBuffer.scala 55:24]
    end else if (io_recv_done) begin // @[IfmBuffer.scala 56:17]
      col_cnt <= 10'h0;
    end else if (io_bram_en_write) begin // @[IfmBuffer.scala 56:38]
      if (col_cnt == _col_cnt_T_1) begin // @[IfmBuffer.scala 56:59]
        col_cnt <= 10'h0;
      end else begin
        col_cnt <= _col_cnt_T_4;
      end
    end
    bram_write_addr_singal <= _GEN_0[10:0]; // @[IfmBuffer.scala 62:{40,40} 64:27]
    bram_write_addr_double <= _GEN_1[10:0]; // @[IfmBuffer.scala 63:{41,41} 65:27]
    temp_single_regnext_0_REG <= temp_single_0[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_0_REG <= temp_double_0[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_1_REG <= temp_single_1[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_1_REG <= temp_double_1[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_2_REG <= temp_single_2[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_2_REG <= temp_double_2[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_3_REG <= temp_single_3[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_3_REG <= temp_double_3[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_4_REG <= temp_single_4[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_4_REG <= temp_double_4[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_5_REG <= temp_single_5[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_5_REG <= temp_double_5[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_6_REG <= temp_single_6[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_6_REG <= temp_double_6[15:8]; // @[IfmBuffer.scala 85:55]
    temp_single_regnext_7_REG <= temp_single_7[15:8]; // @[IfmBuffer.scala 84:55]
    temp_double_regnext_7_REG <= temp_double_7[15:8]; // @[IfmBuffer.scala 85:55]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  in_temp_sel = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  in_temp_0 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  in_temp_1 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  in_temp_2 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  in_temp_3 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  in_temp_4 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  in_temp_5 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  in_temp_6 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  in_temp_7 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  row_is_singal_or_double = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  col_cnt = _RAND_10[9:0];
  _RAND_11 = {1{`RANDOM}};
  bram_write_addr_singal = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  bram_write_addr_double = _RAND_12[10:0];
  _RAND_13 = {1{`RANDOM}};
  temp_single_regnext_0_REG = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  temp_double_regnext_0_REG = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  temp_single_regnext_1_REG = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  temp_double_regnext_1_REG = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  temp_single_regnext_2_REG = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  temp_double_regnext_2_REG = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  temp_single_regnext_3_REG = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  temp_double_regnext_3_REG = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  temp_single_regnext_4_REG = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  temp_double_regnext_4_REG = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  temp_single_regnext_5_REG = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  temp_double_regnext_5_REG = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  temp_single_regnext_6_REG = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  temp_double_regnext_6_REG = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  temp_single_regnext_7_REG = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  temp_double_regnext_7_REG = _RAND_28[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TPRAM_WRAP_16(
  input         clock,
  input         io_wen,
  input  [6:0]  io_waddr,
  input  [6:0]  io_raddr,
  input  [71:0] io_wdata,
  output [71:0] io_rdata
);
  wire  tpram_CLKA; // @[utils.scala 218:23]
  wire  tpram_CLKB; // @[utils.scala 218:23]
  wire  tpram_CENB; // @[utils.scala 218:23]
  wire  tpram_CENA; // @[utils.scala 218:23]
  wire [6:0] tpram_AB; // @[utils.scala 218:23]
  wire [6:0] tpram_AA; // @[utils.scala 218:23]
  wire [71:0] tpram_DB; // @[utils.scala 218:23]
  wire [71:0] tpram_QA; // @[utils.scala 218:23]
  TPRAM #(.DATA_WIDTH(72), .DEPTH(128), .RAM_STYLE_VAL("distributed")) tpram ( // @[utils.scala 218:23]
    .CLKA(tpram_CLKA),
    .CLKB(tpram_CLKB),
    .CENB(tpram_CENB),
    .CENA(tpram_CENA),
    .AB(tpram_AB),
    .AA(tpram_AA),
    .DB(tpram_DB),
    .QA(tpram_QA)
  );
  assign io_rdata = tpram_QA; // @[utils.scala 230:12]
  assign tpram_CLKA = clock; // @[utils.scala 222:19]
  assign tpram_CLKB = clock; // @[utils.scala 223:19]
  assign tpram_CENB = ~io_wen; // @[utils.scala 224:22]
  assign tpram_CENA = 1'h0; // @[utils.scala 225:22]
  assign tpram_AB = io_waddr; // @[utils.scala 226:17]
  assign tpram_AA = io_raddr; // @[utils.scala 227:17]
  assign tpram_DB = io_wdata; // @[utils.scala 228:17]
endmodule
module w_buffer_unit(
  input         clock,
  input  [6:0]  io_write_addr_0,
  input  [6:0]  io_write_addr_1,
  input  [6:0]  io_write_addr_2,
  input  [6:0]  io_write_addr_3,
  input  [6:0]  io_write_addr_4,
  input  [6:0]  io_write_addr_5,
  input  [6:0]  io_write_addr_6,
  input  [6:0]  io_write_addr_7,
  input         io_write_en_0,
  input         io_write_en_1,
  input         io_write_en_2,
  input         io_write_en_3,
  input         io_write_en_4,
  input         io_write_en_5,
  input         io_write_en_6,
  input         io_write_en_7,
  input  [71:0] io_weight_in,
  input  [6:0]  io_read_addr,
  output [71:0] io_weight_out_0,
  output [71:0] io_weight_out_1,
  output [71:0] io_weight_out_2,
  output [71:0] io_weight_out_3,
  output [71:0] io_weight_out_4,
  output [71:0] io_weight_out_5,
  output [71:0] io_weight_out_6,
  output [71:0] io_weight_out_7
);
  wire  TPRAM_WRAP_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_1_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_1_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_1_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_1_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_2_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_2_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_2_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_2_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_3_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_3_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_3_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_3_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_4_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_4_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_4_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_4_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_5_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_5_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_5_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_5_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_6_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_6_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_6_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_6_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_7_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_7_io_raddr; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_7_io_wdata; // @[utils.scala 237:100]
  wire [71:0] TPRAM_WRAP_7_io_rdata; // @[utils.scala 237:100]
  TPRAM_WRAP_16 TPRAM_WRAP ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_clock),
    .io_wen(TPRAM_WRAP_io_wen),
    .io_waddr(TPRAM_WRAP_io_waddr),
    .io_raddr(TPRAM_WRAP_io_raddr),
    .io_wdata(TPRAM_WRAP_io_wdata),
    .io_rdata(TPRAM_WRAP_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_1 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_1_clock),
    .io_wen(TPRAM_WRAP_1_io_wen),
    .io_waddr(TPRAM_WRAP_1_io_waddr),
    .io_raddr(TPRAM_WRAP_1_io_raddr),
    .io_wdata(TPRAM_WRAP_1_io_wdata),
    .io_rdata(TPRAM_WRAP_1_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_2 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_2_clock),
    .io_wen(TPRAM_WRAP_2_io_wen),
    .io_waddr(TPRAM_WRAP_2_io_waddr),
    .io_raddr(TPRAM_WRAP_2_io_raddr),
    .io_wdata(TPRAM_WRAP_2_io_wdata),
    .io_rdata(TPRAM_WRAP_2_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_3 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_3_clock),
    .io_wen(TPRAM_WRAP_3_io_wen),
    .io_waddr(TPRAM_WRAP_3_io_waddr),
    .io_raddr(TPRAM_WRAP_3_io_raddr),
    .io_wdata(TPRAM_WRAP_3_io_wdata),
    .io_rdata(TPRAM_WRAP_3_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_4 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_4_clock),
    .io_wen(TPRAM_WRAP_4_io_wen),
    .io_waddr(TPRAM_WRAP_4_io_waddr),
    .io_raddr(TPRAM_WRAP_4_io_raddr),
    .io_wdata(TPRAM_WRAP_4_io_wdata),
    .io_rdata(TPRAM_WRAP_4_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_5 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_5_clock),
    .io_wen(TPRAM_WRAP_5_io_wen),
    .io_waddr(TPRAM_WRAP_5_io_waddr),
    .io_raddr(TPRAM_WRAP_5_io_raddr),
    .io_wdata(TPRAM_WRAP_5_io_wdata),
    .io_rdata(TPRAM_WRAP_5_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_6 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_6_clock),
    .io_wen(TPRAM_WRAP_6_io_wen),
    .io_waddr(TPRAM_WRAP_6_io_waddr),
    .io_raddr(TPRAM_WRAP_6_io_raddr),
    .io_wdata(TPRAM_WRAP_6_io_wdata),
    .io_rdata(TPRAM_WRAP_6_io_rdata)
  );
  TPRAM_WRAP_16 TPRAM_WRAP_7 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_7_clock),
    .io_wen(TPRAM_WRAP_7_io_wen),
    .io_waddr(TPRAM_WRAP_7_io_waddr),
    .io_raddr(TPRAM_WRAP_7_io_raddr),
    .io_wdata(TPRAM_WRAP_7_io_wdata),
    .io_rdata(TPRAM_WRAP_7_io_rdata)
  );
  assign io_weight_out_0 = TPRAM_WRAP_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_1 = TPRAM_WRAP_1_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_2 = TPRAM_WRAP_2_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_3 = TPRAM_WRAP_3_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_4 = TPRAM_WRAP_4_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_5 = TPRAM_WRAP_5_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_6 = TPRAM_WRAP_6_io_rdata; // @[WeightBuffer.scala 106:26]
  assign io_weight_out_7 = TPRAM_WRAP_7_io_rdata; // @[WeightBuffer.scala 106:26]
  assign TPRAM_WRAP_clock = clock;
  assign TPRAM_WRAP_io_wen = io_write_en_0; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_io_waddr = io_write_addr_0; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_1_clock = clock;
  assign TPRAM_WRAP_1_io_wen = io_write_en_1; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_1_io_waddr = io_write_addr_1; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_1_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_1_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_2_clock = clock;
  assign TPRAM_WRAP_2_io_wen = io_write_en_2; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_2_io_waddr = io_write_addr_2; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_2_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_2_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_3_clock = clock;
  assign TPRAM_WRAP_3_io_wen = io_write_en_3; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_3_io_waddr = io_write_addr_3; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_3_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_3_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_4_clock = clock;
  assign TPRAM_WRAP_4_io_wen = io_write_en_4; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_4_io_waddr = io_write_addr_4; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_4_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_4_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_5_clock = clock;
  assign TPRAM_WRAP_5_io_wen = io_write_en_5; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_5_io_waddr = io_write_addr_5; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_5_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_5_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_6_clock = clock;
  assign TPRAM_WRAP_6_io_wen = io_write_en_6; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_6_io_waddr = io_write_addr_6; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_6_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_6_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
  assign TPRAM_WRAP_7_clock = clock;
  assign TPRAM_WRAP_7_io_wen = io_write_en_7; // @[WeightBuffer.scala 101:20]
  assign TPRAM_WRAP_7_io_waddr = io_write_addr_7; // @[WeightBuffer.scala 103:22]
  assign TPRAM_WRAP_7_io_raddr = io_read_addr; // @[WeightBuffer.scala 104:22]
  assign TPRAM_WRAP_7_io_wdata = io_weight_in; // @[WeightBuffer.scala 105:22]
endmodule
module WeightBuffer(
  input         clock,
  input         reset,
  input         io_clear,
  input         io_bram_write_en,
  input  [7:0]  io_in_0,
  input  [7:0]  io_in_1,
  input  [7:0]  io_in_2,
  input  [7:0]  io_in_3,
  input  [7:0]  io_in_4,
  input  [7:0]  io_in_5,
  input  [7:0]  io_in_6,
  input  [7:0]  io_in_7,
  input  [6:0]  io_read_addr,
  input  [2:0]  io_sel_when_kernal_is_1,
  output [71:0] io_weight_out_0,
  output [71:0] io_weight_out_1,
  output [71:0] io_weight_out_2,
  output [71:0] io_weight_out_3,
  output [71:0] io_weight_out_4,
  output [71:0] io_weight_out_5,
  output [71:0] io_weight_out_6,
  output [71:0] io_weight_out_7,
  output [71:0] io_weight_out_8,
  output [71:0] io_weight_out_9,
  output [71:0] io_weight_out_10,
  output [71:0] io_weight_out_11,
  output [71:0] io_weight_out_12,
  output [71:0] io_weight_out_13,
  output [71:0] io_weight_out_14,
  output [71:0] io_weight_out_15,
  output [71:0] io_weight_out_16,
  output [71:0] io_weight_out_17,
  output [71:0] io_weight_out_18,
  output [71:0] io_weight_out_19,
  output [71:0] io_weight_out_20,
  output [71:0] io_weight_out_21,
  output [71:0] io_weight_out_22,
  output [71:0] io_weight_out_23,
  output [71:0] io_weight_out_24,
  output [71:0] io_weight_out_25,
  output [71:0] io_weight_out_26,
  output [71:0] io_weight_out_27,
  output [71:0] io_weight_out_28,
  output [71:0] io_weight_out_29,
  output [71:0] io_weight_out_30,
  output [71:0] io_weight_out_31,
  output [71:0] io_weight_out_32,
  output [71:0] io_weight_out_33,
  output [71:0] io_weight_out_34,
  output [71:0] io_weight_out_35,
  output [71:0] io_weight_out_36,
  output [71:0] io_weight_out_37,
  output [71:0] io_weight_out_38,
  output [71:0] io_weight_out_39,
  output [71:0] io_weight_out_40,
  output [71:0] io_weight_out_41,
  output [71:0] io_weight_out_42,
  output [71:0] io_weight_out_43,
  output [71:0] io_weight_out_44,
  output [71:0] io_weight_out_45,
  output [71:0] io_weight_out_46,
  output [71:0] io_weight_out_47,
  output [71:0] io_weight_out_48,
  output [71:0] io_weight_out_49,
  output [71:0] io_weight_out_50,
  output [71:0] io_weight_out_51,
  output [71:0] io_weight_out_52,
  output [71:0] io_weight_out_53,
  output [71:0] io_weight_out_54,
  output [71:0] io_weight_out_55,
  output [71:0] io_weight_out_56,
  output [71:0] io_weight_out_57,
  output [71:0] io_weight_out_58,
  output [71:0] io_weight_out_59,
  output [71:0] io_weight_out_60,
  output [71:0] io_weight_out_61,
  output [71:0] io_weight_out_62,
  output [71:0] io_weight_out_63,
  input         io_kernal
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
`endif // RANDOMIZE_REG_INIT
  wire  buf_unit_0_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_0_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_0_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_0_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_1_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_1_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_1_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_2_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_2_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_2_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_3_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_3_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_3_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_4_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_4_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_4_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_5_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_5_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_5_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_6_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_6_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_6_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_clock; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_0; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_1; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_2; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_3; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_4; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_5; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_6; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_write_addr_7; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_0; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_1; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_2; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_3; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_4; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_5; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_6; // @[WeightBuffer.scala 76:42]
  wire  buf_unit_7_io_write_en_7; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_in; // @[WeightBuffer.scala 76:42]
  wire [6:0] buf_unit_7_io_read_addr; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_0; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_1; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_2; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_3; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_4; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_5; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_6; // @[WeightBuffer.scala 76:42]
  wire [71:0] buf_unit_7_io_weight_out_7; // @[WeightBuffer.scala 76:42]
  reg [7:0] temp_0_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_0_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_1_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_2_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_3_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_4_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_5_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_6_8; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_0; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_1; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_2; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_3; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_4; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_5; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_6; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_7; // @[WeightBuffer.scala 17:51]
  reg [7:0] temp_7_8; // @[WeightBuffer.scala 17:51]
  wire [71:0] w_data_when_k_is_3_0 = {temp_0_0,temp_0_1,temp_0_2,temp_0_3,temp_0_4,temp_0_5,temp_0_6,temp_0_7,temp_0_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_0 = {8'h0,w_data_when_k_is_3_0[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_1 = {temp_1_0,temp_1_1,temp_1_2,temp_1_3,temp_1_4,temp_1_5,temp_1_6,temp_1_7,temp_1_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_1 = {8'h0,w_data_when_k_is_3_1[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_2 = {temp_2_0,temp_2_1,temp_2_2,temp_2_3,temp_2_4,temp_2_5,temp_2_6,temp_2_7,temp_2_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_2 = {8'h0,w_data_when_k_is_3_2[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_3 = {temp_3_0,temp_3_1,temp_3_2,temp_3_3,temp_3_4,temp_3_5,temp_3_6,temp_3_7,temp_3_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_3 = {8'h0,w_data_when_k_is_3_3[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_4 = {temp_4_0,temp_4_1,temp_4_2,temp_4_3,temp_4_4,temp_4_5,temp_4_6,temp_4_7,temp_4_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_4 = {8'h0,w_data_when_k_is_3_4[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_5 = {temp_5_0,temp_5_1,temp_5_2,temp_5_3,temp_5_4,temp_5_5,temp_5_6,temp_5_7,temp_5_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_5 = {8'h0,w_data_when_k_is_3_5[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_6 = {temp_6_0,temp_6_1,temp_6_2,temp_6_3,temp_6_4,temp_6_5,temp_6_6,temp_6_7,temp_6_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_6 = {8'h0,w_data_when_k_is_3_6[63:0]}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_3_7 = {temp_7_0,temp_7_1,temp_7_2,temp_7_3,temp_7_4,temp_7_5,temp_7_6,temp_7_7,temp_7_8}; // @[Cat.scala 33:92]
  wire [71:0] w_data_when_k_is_1_7 = {8'h0,w_data_when_k_is_3_7[63:0]}; // @[Cat.scala 33:92]
  reg [3:0] cnt9; // @[WeightBuffer.scala 42:23]
  wire [3:0] cnt9_max = io_kernal ? 4'h8 : 4'h7; // @[WeightBuffer.scala 43:23]
  reg [2:0] cnt8; // @[WeightBuffer.scala 44:23]
  wire  rst = reset | io_clear; // @[WeightBuffer.scala 45:28]
  wire  _cnt9_T = cnt9 == cnt9_max; // @[WeightBuffer.scala 46:58]
  wire [3:0] _cnt9_T_2 = cnt9 + 4'h1; // @[WeightBuffer.scala 46:82]
  wire  _cnt8_T_1 = cnt8 == 3'h7; // @[WeightBuffer.scala 47:83]
  wire [2:0] _cnt8_T_3 = cnt8 + 3'h1; // @[WeightBuffer.scala 47:111]
  wire [2:0] _cnt8_T_4 = cnt8 == 3'h7 ? 3'h0 : _cnt8_T_3; // @[WeightBuffer.scala 47:77]
  reg  ch_en_reg_0; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_1; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_2; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_3; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_4; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_5; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_6; // @[WeightBuffer.scala 49:24]
  reg  ch_en_reg_7; // @[WeightBuffer.scala 49:24]
  wire  _ch_en_0_T = cnt8 == 3'h0; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_1_T = cnt8 == 3'h1; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_2_T = cnt8 == 3'h2; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_3_T = cnt8 == 3'h3; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_4_T = cnt8 == 3'h4; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_5_T = cnt8 == 3'h5; // @[WeightBuffer.scala 51:47]
  wire  _ch_en_6_T = cnt8 == 3'h6; // @[WeightBuffer.scala 51:47]
  reg [6:0] ch_cnt_0; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_1; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_2; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_3; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_4; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_5; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_6; // @[WeightBuffer.scala 55:40]
  reg [6:0] ch_cnt_7; // @[WeightBuffer.scala 55:40]
  wire [6:0] _ch_cnt_0_T_1 = ch_cnt_0 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_1_T_1 = ch_cnt_1 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_2_T_1 = ch_cnt_2 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_3_T_1 = ch_cnt_3 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_4_T_1 = ch_cnt_4 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_5_T_1 = ch_cnt_5 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_6_T_1 = ch_cnt_6 + 7'h1; // @[WeightBuffer.scala 57:64]
  wire [6:0] _ch_cnt_7_T_1 = ch_cnt_7 + 7'h1; // @[WeightBuffer.scala 57:64]
  reg  bram_write_en_downedge_REG; // @[utils.scala 19:16]
  wire  bram_write_en_downedge = bram_write_en_downedge_REG & ~io_bram_write_en; // @[utils.scala 19:26]
  wire  force_write_0 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_0_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_1 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_1_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_2 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_2_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_3 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_3_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_4 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_4_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_5 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_5_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_6 = bram_write_en_downedge & cnt9 != 4'h0 & _ch_en_6_T; // @[WeightBuffer.scala 63:61]
  wire  force_write_7 = bram_write_en_downedge & cnt9 != 4'h0 & _cnt8_T_1; // @[WeightBuffer.scala 63:61]
  wire [71:0] weight_out_0 = buf_unit_0_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_0_0 = weight_out_0[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_1 = weight_out_0[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_2 = weight_out_0[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_3 = weight_out_0[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_4 = weight_out_0[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_5 = weight_out_0[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_6 = weight_out_0[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_0_7 = weight_out_0[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_73 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_0_1 : read_data_0_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_74 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_0_2 : _GEN_73; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_75 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_0_3 : _GEN_74; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_76 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_0_4 : _GEN_75; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_77 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_0_5 : _GEN_76; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_78 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_0_6 : _GEN_77; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_0 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_0_7 : _GEN_78; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_1 = buf_unit_0_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_1_0 = weight_out_1[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_1 = weight_out_1[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_2 = weight_out_1[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_3 = weight_out_1[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_4 = weight_out_1[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_5 = weight_out_1[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_6 = weight_out_1[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_1_7 = weight_out_1[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_81 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_1_1 : read_data_1_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_82 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_1_2 : _GEN_81; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_83 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_1_3 : _GEN_82; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_84 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_1_4 : _GEN_83; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_85 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_1_5 : _GEN_84; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_86 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_1_6 : _GEN_85; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_1 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_1_7 : _GEN_86; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_2 = buf_unit_0_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_2_0 = weight_out_2[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_1 = weight_out_2[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_2 = weight_out_2[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_3 = weight_out_2[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_4 = weight_out_2[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_5 = weight_out_2[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_6 = weight_out_2[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_2_7 = weight_out_2[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_89 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_2_1 : read_data_2_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_90 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_2_2 : _GEN_89; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_91 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_2_3 : _GEN_90; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_92 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_2_4 : _GEN_91; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_93 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_2_5 : _GEN_92; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_94 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_2_6 : _GEN_93; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_2 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_2_7 : _GEN_94; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_3 = buf_unit_0_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_3_0 = weight_out_3[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_1 = weight_out_3[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_2 = weight_out_3[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_3 = weight_out_3[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_4 = weight_out_3[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_5 = weight_out_3[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_6 = weight_out_3[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_3_7 = weight_out_3[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_97 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_3_1 : read_data_3_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_98 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_3_2 : _GEN_97; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_99 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_3_3 : _GEN_98; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_100 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_3_4 : _GEN_99; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_101 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_3_5 : _GEN_100; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_102 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_3_6 : _GEN_101; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_3 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_3_7 : _GEN_102; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_4 = buf_unit_0_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_4_0 = weight_out_4[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_1 = weight_out_4[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_2 = weight_out_4[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_3 = weight_out_4[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_4 = weight_out_4[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_5 = weight_out_4[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_6 = weight_out_4[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_4_7 = weight_out_4[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_105 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_4_1 : read_data_4_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_106 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_4_2 : _GEN_105; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_107 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_4_3 : _GEN_106; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_108 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_4_4 : _GEN_107; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_109 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_4_5 : _GEN_108; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_110 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_4_6 : _GEN_109; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_4 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_4_7 : _GEN_110; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_5 = buf_unit_0_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_5_0 = weight_out_5[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_1 = weight_out_5[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_2 = weight_out_5[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_3 = weight_out_5[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_4 = weight_out_5[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_5 = weight_out_5[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_6 = weight_out_5[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_5_7 = weight_out_5[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_113 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_5_1 : read_data_5_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_114 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_5_2 : _GEN_113; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_115 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_5_3 : _GEN_114; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_116 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_5_4 : _GEN_115; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_117 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_5_5 : _GEN_116; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_118 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_5_6 : _GEN_117; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_5 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_5_7 : _GEN_118; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_6 = buf_unit_0_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_6_0 = weight_out_6[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_1 = weight_out_6[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_2 = weight_out_6[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_3 = weight_out_6[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_4 = weight_out_6[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_5 = weight_out_6[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_6 = weight_out_6[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_6_7 = weight_out_6[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_121 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_6_1 : read_data_6_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_122 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_6_2 : _GEN_121; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_123 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_6_3 : _GEN_122; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_124 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_6_4 : _GEN_123; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_125 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_6_5 : _GEN_124; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_126 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_6_6 : _GEN_125; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_6 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_6_7 : _GEN_126; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_7 = buf_unit_0_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_7_0 = weight_out_7[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_1 = weight_out_7[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_2 = weight_out_7[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_3 = weight_out_7[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_4 = weight_out_7[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_5 = weight_out_7[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_6 = weight_out_7[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_7_7 = weight_out_7[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_129 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_7_1 : read_data_7_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_130 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_7_2 : _GEN_129; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_131 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_7_3 : _GEN_130; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_132 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_7_4 : _GEN_131; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_133 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_7_5 : _GEN_132; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_134 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_7_6 : _GEN_133; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_7 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_7_7 : _GEN_134; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_8 = buf_unit_1_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_8_0 = weight_out_8[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_1 = weight_out_8[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_2 = weight_out_8[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_3 = weight_out_8[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_4 = weight_out_8[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_5 = weight_out_8[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_6 = weight_out_8[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_8_7 = weight_out_8[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_137 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_8_1 : read_data_8_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_138 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_8_2 : _GEN_137; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_139 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_8_3 : _GEN_138; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_140 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_8_4 : _GEN_139; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_141 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_8_5 : _GEN_140; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_142 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_8_6 : _GEN_141; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_8 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_8_7 : _GEN_142; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_9 = buf_unit_1_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_9_0 = weight_out_9[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_1 = weight_out_9[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_2 = weight_out_9[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_3 = weight_out_9[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_4 = weight_out_9[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_5 = weight_out_9[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_6 = weight_out_9[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_9_7 = weight_out_9[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_145 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_9_1 : read_data_9_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_146 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_9_2 : _GEN_145; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_147 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_9_3 : _GEN_146; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_148 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_9_4 : _GEN_147; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_149 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_9_5 : _GEN_148; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_150 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_9_6 : _GEN_149; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_9 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_9_7 : _GEN_150; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_10 = buf_unit_1_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_10_0 = weight_out_10[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_1 = weight_out_10[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_2 = weight_out_10[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_3 = weight_out_10[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_4 = weight_out_10[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_5 = weight_out_10[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_6 = weight_out_10[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_10_7 = weight_out_10[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_153 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_10_1 : read_data_10_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_154 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_10_2 : _GEN_153; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_155 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_10_3 : _GEN_154; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_156 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_10_4 : _GEN_155; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_157 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_10_5 : _GEN_156; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_158 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_10_6 : _GEN_157; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_10 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_10_7 : _GEN_158; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_11 = buf_unit_1_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_11_0 = weight_out_11[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_1 = weight_out_11[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_2 = weight_out_11[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_3 = weight_out_11[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_4 = weight_out_11[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_5 = weight_out_11[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_6 = weight_out_11[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_11_7 = weight_out_11[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_161 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_11_1 : read_data_11_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_162 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_11_2 : _GEN_161; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_163 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_11_3 : _GEN_162; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_164 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_11_4 : _GEN_163; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_165 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_11_5 : _GEN_164; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_166 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_11_6 : _GEN_165; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_11 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_11_7 : _GEN_166; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_12 = buf_unit_1_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_12_0 = weight_out_12[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_1 = weight_out_12[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_2 = weight_out_12[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_3 = weight_out_12[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_4 = weight_out_12[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_5 = weight_out_12[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_6 = weight_out_12[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_12_7 = weight_out_12[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_169 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_12_1 : read_data_12_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_170 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_12_2 : _GEN_169; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_171 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_12_3 : _GEN_170; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_172 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_12_4 : _GEN_171; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_173 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_12_5 : _GEN_172; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_174 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_12_6 : _GEN_173; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_12 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_12_7 : _GEN_174; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_13 = buf_unit_1_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_13_0 = weight_out_13[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_1 = weight_out_13[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_2 = weight_out_13[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_3 = weight_out_13[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_4 = weight_out_13[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_5 = weight_out_13[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_6 = weight_out_13[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_13_7 = weight_out_13[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_177 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_13_1 : read_data_13_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_178 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_13_2 : _GEN_177; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_179 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_13_3 : _GEN_178; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_180 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_13_4 : _GEN_179; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_181 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_13_5 : _GEN_180; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_182 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_13_6 : _GEN_181; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_13 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_13_7 : _GEN_182; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_14 = buf_unit_1_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_14_0 = weight_out_14[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_1 = weight_out_14[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_2 = weight_out_14[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_3 = weight_out_14[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_4 = weight_out_14[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_5 = weight_out_14[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_6 = weight_out_14[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_14_7 = weight_out_14[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_185 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_14_1 : read_data_14_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_186 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_14_2 : _GEN_185; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_187 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_14_3 : _GEN_186; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_188 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_14_4 : _GEN_187; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_189 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_14_5 : _GEN_188; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_190 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_14_6 : _GEN_189; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_14 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_14_7 : _GEN_190; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_15 = buf_unit_1_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_15_0 = weight_out_15[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_1 = weight_out_15[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_2 = weight_out_15[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_3 = weight_out_15[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_4 = weight_out_15[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_5 = weight_out_15[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_6 = weight_out_15[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_15_7 = weight_out_15[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_193 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_15_1 : read_data_15_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_194 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_15_2 : _GEN_193; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_195 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_15_3 : _GEN_194; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_196 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_15_4 : _GEN_195; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_197 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_15_5 : _GEN_196; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_198 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_15_6 : _GEN_197; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_15 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_15_7 : _GEN_198; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_16 = buf_unit_2_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_16_0 = weight_out_16[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_1 = weight_out_16[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_2 = weight_out_16[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_3 = weight_out_16[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_4 = weight_out_16[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_5 = weight_out_16[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_6 = weight_out_16[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_16_7 = weight_out_16[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_201 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_16_1 : read_data_16_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_202 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_16_2 : _GEN_201; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_203 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_16_3 : _GEN_202; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_204 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_16_4 : _GEN_203; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_205 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_16_5 : _GEN_204; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_206 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_16_6 : _GEN_205; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_16 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_16_7 : _GEN_206; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_17 = buf_unit_2_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_17_0 = weight_out_17[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_1 = weight_out_17[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_2 = weight_out_17[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_3 = weight_out_17[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_4 = weight_out_17[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_5 = weight_out_17[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_6 = weight_out_17[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_17_7 = weight_out_17[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_209 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_17_1 : read_data_17_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_210 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_17_2 : _GEN_209; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_211 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_17_3 : _GEN_210; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_212 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_17_4 : _GEN_211; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_213 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_17_5 : _GEN_212; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_214 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_17_6 : _GEN_213; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_17 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_17_7 : _GEN_214; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_18 = buf_unit_2_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_18_0 = weight_out_18[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_1 = weight_out_18[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_2 = weight_out_18[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_3 = weight_out_18[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_4 = weight_out_18[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_5 = weight_out_18[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_6 = weight_out_18[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_18_7 = weight_out_18[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_217 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_18_1 : read_data_18_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_218 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_18_2 : _GEN_217; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_219 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_18_3 : _GEN_218; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_220 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_18_4 : _GEN_219; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_221 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_18_5 : _GEN_220; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_222 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_18_6 : _GEN_221; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_18 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_18_7 : _GEN_222; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_19 = buf_unit_2_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_19_0 = weight_out_19[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_1 = weight_out_19[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_2 = weight_out_19[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_3 = weight_out_19[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_4 = weight_out_19[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_5 = weight_out_19[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_6 = weight_out_19[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_19_7 = weight_out_19[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_225 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_19_1 : read_data_19_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_226 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_19_2 : _GEN_225; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_227 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_19_3 : _GEN_226; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_228 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_19_4 : _GEN_227; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_229 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_19_5 : _GEN_228; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_230 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_19_6 : _GEN_229; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_19 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_19_7 : _GEN_230; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_20 = buf_unit_2_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_20_0 = weight_out_20[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_1 = weight_out_20[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_2 = weight_out_20[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_3 = weight_out_20[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_4 = weight_out_20[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_5 = weight_out_20[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_6 = weight_out_20[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_20_7 = weight_out_20[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_233 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_20_1 : read_data_20_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_234 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_20_2 : _GEN_233; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_235 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_20_3 : _GEN_234; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_236 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_20_4 : _GEN_235; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_237 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_20_5 : _GEN_236; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_238 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_20_6 : _GEN_237; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_20 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_20_7 : _GEN_238; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_21 = buf_unit_2_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_21_0 = weight_out_21[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_1 = weight_out_21[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_2 = weight_out_21[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_3 = weight_out_21[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_4 = weight_out_21[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_5 = weight_out_21[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_6 = weight_out_21[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_21_7 = weight_out_21[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_241 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_21_1 : read_data_21_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_242 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_21_2 : _GEN_241; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_243 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_21_3 : _GEN_242; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_244 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_21_4 : _GEN_243; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_245 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_21_5 : _GEN_244; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_246 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_21_6 : _GEN_245; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_21 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_21_7 : _GEN_246; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_22 = buf_unit_2_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_22_0 = weight_out_22[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_1 = weight_out_22[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_2 = weight_out_22[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_3 = weight_out_22[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_4 = weight_out_22[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_5 = weight_out_22[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_6 = weight_out_22[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_22_7 = weight_out_22[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_249 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_22_1 : read_data_22_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_250 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_22_2 : _GEN_249; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_251 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_22_3 : _GEN_250; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_252 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_22_4 : _GEN_251; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_253 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_22_5 : _GEN_252; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_254 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_22_6 : _GEN_253; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_22 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_22_7 : _GEN_254; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_23 = buf_unit_2_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_23_0 = weight_out_23[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_1 = weight_out_23[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_2 = weight_out_23[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_3 = weight_out_23[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_4 = weight_out_23[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_5 = weight_out_23[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_6 = weight_out_23[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_23_7 = weight_out_23[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_257 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_23_1 : read_data_23_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_258 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_23_2 : _GEN_257; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_259 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_23_3 : _GEN_258; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_260 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_23_4 : _GEN_259; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_261 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_23_5 : _GEN_260; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_262 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_23_6 : _GEN_261; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_23 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_23_7 : _GEN_262; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_24 = buf_unit_3_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_24_0 = weight_out_24[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_1 = weight_out_24[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_2 = weight_out_24[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_3 = weight_out_24[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_4 = weight_out_24[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_5 = weight_out_24[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_6 = weight_out_24[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_24_7 = weight_out_24[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_265 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_24_1 : read_data_24_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_266 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_24_2 : _GEN_265; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_267 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_24_3 : _GEN_266; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_268 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_24_4 : _GEN_267; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_269 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_24_5 : _GEN_268; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_270 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_24_6 : _GEN_269; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_24 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_24_7 : _GEN_270; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_25 = buf_unit_3_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_25_0 = weight_out_25[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_1 = weight_out_25[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_2 = weight_out_25[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_3 = weight_out_25[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_4 = weight_out_25[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_5 = weight_out_25[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_6 = weight_out_25[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_25_7 = weight_out_25[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_273 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_25_1 : read_data_25_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_274 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_25_2 : _GEN_273; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_275 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_25_3 : _GEN_274; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_276 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_25_4 : _GEN_275; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_277 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_25_5 : _GEN_276; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_278 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_25_6 : _GEN_277; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_25 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_25_7 : _GEN_278; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_26 = buf_unit_3_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_26_0 = weight_out_26[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_1 = weight_out_26[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_2 = weight_out_26[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_3 = weight_out_26[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_4 = weight_out_26[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_5 = weight_out_26[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_6 = weight_out_26[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_26_7 = weight_out_26[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_281 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_26_1 : read_data_26_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_282 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_26_2 : _GEN_281; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_283 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_26_3 : _GEN_282; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_284 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_26_4 : _GEN_283; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_285 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_26_5 : _GEN_284; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_286 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_26_6 : _GEN_285; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_26 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_26_7 : _GEN_286; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_27 = buf_unit_3_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_27_0 = weight_out_27[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_1 = weight_out_27[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_2 = weight_out_27[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_3 = weight_out_27[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_4 = weight_out_27[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_5 = weight_out_27[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_6 = weight_out_27[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_27_7 = weight_out_27[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_289 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_27_1 : read_data_27_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_290 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_27_2 : _GEN_289; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_291 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_27_3 : _GEN_290; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_292 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_27_4 : _GEN_291; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_293 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_27_5 : _GEN_292; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_294 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_27_6 : _GEN_293; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_27 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_27_7 : _GEN_294; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_28 = buf_unit_3_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_28_0 = weight_out_28[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_1 = weight_out_28[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_2 = weight_out_28[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_3 = weight_out_28[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_4 = weight_out_28[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_5 = weight_out_28[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_6 = weight_out_28[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_28_7 = weight_out_28[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_297 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_28_1 : read_data_28_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_298 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_28_2 : _GEN_297; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_299 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_28_3 : _GEN_298; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_300 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_28_4 : _GEN_299; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_301 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_28_5 : _GEN_300; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_302 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_28_6 : _GEN_301; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_28 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_28_7 : _GEN_302; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_29 = buf_unit_3_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_29_0 = weight_out_29[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_1 = weight_out_29[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_2 = weight_out_29[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_3 = weight_out_29[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_4 = weight_out_29[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_5 = weight_out_29[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_6 = weight_out_29[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_29_7 = weight_out_29[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_305 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_29_1 : read_data_29_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_306 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_29_2 : _GEN_305; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_307 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_29_3 : _GEN_306; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_308 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_29_4 : _GEN_307; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_309 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_29_5 : _GEN_308; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_310 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_29_6 : _GEN_309; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_29 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_29_7 : _GEN_310; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_30 = buf_unit_3_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_30_0 = weight_out_30[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_1 = weight_out_30[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_2 = weight_out_30[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_3 = weight_out_30[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_4 = weight_out_30[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_5 = weight_out_30[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_6 = weight_out_30[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_30_7 = weight_out_30[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_313 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_30_1 : read_data_30_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_314 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_30_2 : _GEN_313; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_315 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_30_3 : _GEN_314; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_316 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_30_4 : _GEN_315; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_317 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_30_5 : _GEN_316; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_318 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_30_6 : _GEN_317; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_30 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_30_7 : _GEN_318; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_31 = buf_unit_3_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_31_0 = weight_out_31[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_1 = weight_out_31[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_2 = weight_out_31[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_3 = weight_out_31[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_4 = weight_out_31[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_5 = weight_out_31[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_6 = weight_out_31[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_31_7 = weight_out_31[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_321 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_31_1 : read_data_31_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_322 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_31_2 : _GEN_321; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_323 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_31_3 : _GEN_322; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_324 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_31_4 : _GEN_323; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_325 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_31_5 : _GEN_324; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_326 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_31_6 : _GEN_325; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_31 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_31_7 : _GEN_326; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_32 = buf_unit_4_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_32_0 = weight_out_32[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_1 = weight_out_32[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_2 = weight_out_32[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_3 = weight_out_32[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_4 = weight_out_32[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_5 = weight_out_32[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_6 = weight_out_32[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_32_7 = weight_out_32[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_329 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_32_1 : read_data_32_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_330 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_32_2 : _GEN_329; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_331 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_32_3 : _GEN_330; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_332 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_32_4 : _GEN_331; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_333 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_32_5 : _GEN_332; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_334 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_32_6 : _GEN_333; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_32 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_32_7 : _GEN_334; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_33 = buf_unit_4_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_33_0 = weight_out_33[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_1 = weight_out_33[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_2 = weight_out_33[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_3 = weight_out_33[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_4 = weight_out_33[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_5 = weight_out_33[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_6 = weight_out_33[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_33_7 = weight_out_33[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_337 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_33_1 : read_data_33_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_338 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_33_2 : _GEN_337; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_339 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_33_3 : _GEN_338; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_340 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_33_4 : _GEN_339; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_341 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_33_5 : _GEN_340; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_342 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_33_6 : _GEN_341; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_33 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_33_7 : _GEN_342; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_34 = buf_unit_4_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_34_0 = weight_out_34[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_1 = weight_out_34[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_2 = weight_out_34[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_3 = weight_out_34[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_4 = weight_out_34[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_5 = weight_out_34[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_6 = weight_out_34[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_34_7 = weight_out_34[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_345 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_34_1 : read_data_34_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_346 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_34_2 : _GEN_345; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_347 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_34_3 : _GEN_346; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_348 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_34_4 : _GEN_347; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_349 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_34_5 : _GEN_348; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_350 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_34_6 : _GEN_349; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_34 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_34_7 : _GEN_350; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_35 = buf_unit_4_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_35_0 = weight_out_35[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_1 = weight_out_35[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_2 = weight_out_35[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_3 = weight_out_35[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_4 = weight_out_35[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_5 = weight_out_35[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_6 = weight_out_35[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_35_7 = weight_out_35[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_353 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_35_1 : read_data_35_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_354 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_35_2 : _GEN_353; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_355 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_35_3 : _GEN_354; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_356 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_35_4 : _GEN_355; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_357 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_35_5 : _GEN_356; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_358 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_35_6 : _GEN_357; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_35 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_35_7 : _GEN_358; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_36 = buf_unit_4_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_36_0 = weight_out_36[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_1 = weight_out_36[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_2 = weight_out_36[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_3 = weight_out_36[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_4 = weight_out_36[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_5 = weight_out_36[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_6 = weight_out_36[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_36_7 = weight_out_36[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_361 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_36_1 : read_data_36_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_362 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_36_2 : _GEN_361; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_363 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_36_3 : _GEN_362; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_364 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_36_4 : _GEN_363; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_365 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_36_5 : _GEN_364; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_366 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_36_6 : _GEN_365; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_36 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_36_7 : _GEN_366; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_37 = buf_unit_4_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_37_0 = weight_out_37[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_1 = weight_out_37[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_2 = weight_out_37[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_3 = weight_out_37[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_4 = weight_out_37[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_5 = weight_out_37[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_6 = weight_out_37[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_37_7 = weight_out_37[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_369 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_37_1 : read_data_37_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_370 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_37_2 : _GEN_369; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_371 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_37_3 : _GEN_370; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_372 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_37_4 : _GEN_371; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_373 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_37_5 : _GEN_372; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_374 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_37_6 : _GEN_373; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_37 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_37_7 : _GEN_374; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_38 = buf_unit_4_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_38_0 = weight_out_38[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_1 = weight_out_38[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_2 = weight_out_38[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_3 = weight_out_38[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_4 = weight_out_38[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_5 = weight_out_38[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_6 = weight_out_38[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_38_7 = weight_out_38[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_377 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_38_1 : read_data_38_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_378 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_38_2 : _GEN_377; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_379 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_38_3 : _GEN_378; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_380 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_38_4 : _GEN_379; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_381 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_38_5 : _GEN_380; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_382 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_38_6 : _GEN_381; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_38 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_38_7 : _GEN_382; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_39 = buf_unit_4_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_39_0 = weight_out_39[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_1 = weight_out_39[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_2 = weight_out_39[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_3 = weight_out_39[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_4 = weight_out_39[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_5 = weight_out_39[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_6 = weight_out_39[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_39_7 = weight_out_39[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_385 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_39_1 : read_data_39_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_386 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_39_2 : _GEN_385; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_387 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_39_3 : _GEN_386; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_388 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_39_4 : _GEN_387; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_389 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_39_5 : _GEN_388; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_390 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_39_6 : _GEN_389; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_39 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_39_7 : _GEN_390; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_40 = buf_unit_5_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_40_0 = weight_out_40[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_1 = weight_out_40[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_2 = weight_out_40[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_3 = weight_out_40[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_4 = weight_out_40[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_5 = weight_out_40[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_6 = weight_out_40[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_40_7 = weight_out_40[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_393 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_40_1 : read_data_40_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_394 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_40_2 : _GEN_393; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_395 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_40_3 : _GEN_394; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_396 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_40_4 : _GEN_395; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_397 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_40_5 : _GEN_396; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_398 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_40_6 : _GEN_397; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_40 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_40_7 : _GEN_398; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_41 = buf_unit_5_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_41_0 = weight_out_41[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_1 = weight_out_41[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_2 = weight_out_41[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_3 = weight_out_41[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_4 = weight_out_41[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_5 = weight_out_41[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_6 = weight_out_41[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_41_7 = weight_out_41[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_401 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_41_1 : read_data_41_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_402 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_41_2 : _GEN_401; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_403 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_41_3 : _GEN_402; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_404 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_41_4 : _GEN_403; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_405 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_41_5 : _GEN_404; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_406 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_41_6 : _GEN_405; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_41 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_41_7 : _GEN_406; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_42 = buf_unit_5_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_42_0 = weight_out_42[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_1 = weight_out_42[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_2 = weight_out_42[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_3 = weight_out_42[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_4 = weight_out_42[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_5 = weight_out_42[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_6 = weight_out_42[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_42_7 = weight_out_42[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_409 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_42_1 : read_data_42_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_410 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_42_2 : _GEN_409; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_411 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_42_3 : _GEN_410; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_412 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_42_4 : _GEN_411; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_413 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_42_5 : _GEN_412; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_414 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_42_6 : _GEN_413; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_42 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_42_7 : _GEN_414; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_43 = buf_unit_5_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_43_0 = weight_out_43[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_1 = weight_out_43[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_2 = weight_out_43[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_3 = weight_out_43[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_4 = weight_out_43[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_5 = weight_out_43[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_6 = weight_out_43[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_43_7 = weight_out_43[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_417 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_43_1 : read_data_43_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_418 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_43_2 : _GEN_417; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_419 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_43_3 : _GEN_418; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_420 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_43_4 : _GEN_419; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_421 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_43_5 : _GEN_420; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_422 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_43_6 : _GEN_421; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_43 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_43_7 : _GEN_422; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_44 = buf_unit_5_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_44_0 = weight_out_44[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_1 = weight_out_44[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_2 = weight_out_44[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_3 = weight_out_44[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_4 = weight_out_44[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_5 = weight_out_44[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_6 = weight_out_44[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_44_7 = weight_out_44[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_425 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_44_1 : read_data_44_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_426 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_44_2 : _GEN_425; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_427 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_44_3 : _GEN_426; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_428 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_44_4 : _GEN_427; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_429 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_44_5 : _GEN_428; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_430 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_44_6 : _GEN_429; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_44 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_44_7 : _GEN_430; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_45 = buf_unit_5_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_45_0 = weight_out_45[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_1 = weight_out_45[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_2 = weight_out_45[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_3 = weight_out_45[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_4 = weight_out_45[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_5 = weight_out_45[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_6 = weight_out_45[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_45_7 = weight_out_45[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_433 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_45_1 : read_data_45_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_434 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_45_2 : _GEN_433; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_435 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_45_3 : _GEN_434; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_436 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_45_4 : _GEN_435; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_437 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_45_5 : _GEN_436; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_438 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_45_6 : _GEN_437; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_45 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_45_7 : _GEN_438; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_46 = buf_unit_5_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_46_0 = weight_out_46[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_1 = weight_out_46[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_2 = weight_out_46[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_3 = weight_out_46[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_4 = weight_out_46[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_5 = weight_out_46[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_6 = weight_out_46[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_46_7 = weight_out_46[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_441 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_46_1 : read_data_46_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_442 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_46_2 : _GEN_441; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_443 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_46_3 : _GEN_442; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_444 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_46_4 : _GEN_443; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_445 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_46_5 : _GEN_444; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_446 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_46_6 : _GEN_445; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_46 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_46_7 : _GEN_446; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_47 = buf_unit_5_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_47_0 = weight_out_47[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_1 = weight_out_47[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_2 = weight_out_47[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_3 = weight_out_47[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_4 = weight_out_47[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_5 = weight_out_47[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_6 = weight_out_47[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_47_7 = weight_out_47[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_449 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_47_1 : read_data_47_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_450 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_47_2 : _GEN_449; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_451 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_47_3 : _GEN_450; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_452 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_47_4 : _GEN_451; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_453 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_47_5 : _GEN_452; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_454 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_47_6 : _GEN_453; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_47 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_47_7 : _GEN_454; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_48 = buf_unit_6_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_48_0 = weight_out_48[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_1 = weight_out_48[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_2 = weight_out_48[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_3 = weight_out_48[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_4 = weight_out_48[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_5 = weight_out_48[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_6 = weight_out_48[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_48_7 = weight_out_48[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_457 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_48_1 : read_data_48_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_458 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_48_2 : _GEN_457; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_459 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_48_3 : _GEN_458; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_460 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_48_4 : _GEN_459; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_461 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_48_5 : _GEN_460; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_462 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_48_6 : _GEN_461; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_48 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_48_7 : _GEN_462; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_49 = buf_unit_6_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_49_0 = weight_out_49[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_1 = weight_out_49[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_2 = weight_out_49[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_3 = weight_out_49[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_4 = weight_out_49[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_5 = weight_out_49[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_6 = weight_out_49[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_49_7 = weight_out_49[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_465 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_49_1 : read_data_49_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_466 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_49_2 : _GEN_465; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_467 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_49_3 : _GEN_466; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_468 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_49_4 : _GEN_467; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_469 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_49_5 : _GEN_468; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_470 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_49_6 : _GEN_469; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_49 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_49_7 : _GEN_470; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_50 = buf_unit_6_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_50_0 = weight_out_50[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_1 = weight_out_50[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_2 = weight_out_50[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_3 = weight_out_50[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_4 = weight_out_50[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_5 = weight_out_50[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_6 = weight_out_50[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_50_7 = weight_out_50[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_473 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_50_1 : read_data_50_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_474 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_50_2 : _GEN_473; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_475 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_50_3 : _GEN_474; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_476 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_50_4 : _GEN_475; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_477 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_50_5 : _GEN_476; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_478 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_50_6 : _GEN_477; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_50 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_50_7 : _GEN_478; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_51 = buf_unit_6_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_51_0 = weight_out_51[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_1 = weight_out_51[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_2 = weight_out_51[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_3 = weight_out_51[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_4 = weight_out_51[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_5 = weight_out_51[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_6 = weight_out_51[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_51_7 = weight_out_51[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_481 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_51_1 : read_data_51_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_482 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_51_2 : _GEN_481; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_483 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_51_3 : _GEN_482; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_484 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_51_4 : _GEN_483; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_485 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_51_5 : _GEN_484; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_486 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_51_6 : _GEN_485; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_51 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_51_7 : _GEN_486; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_52 = buf_unit_6_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_52_0 = weight_out_52[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_1 = weight_out_52[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_2 = weight_out_52[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_3 = weight_out_52[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_4 = weight_out_52[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_5 = weight_out_52[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_6 = weight_out_52[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_52_7 = weight_out_52[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_489 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_52_1 : read_data_52_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_490 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_52_2 : _GEN_489; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_491 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_52_3 : _GEN_490; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_492 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_52_4 : _GEN_491; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_493 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_52_5 : _GEN_492; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_494 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_52_6 : _GEN_493; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_52 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_52_7 : _GEN_494; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_53 = buf_unit_6_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_53_0 = weight_out_53[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_1 = weight_out_53[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_2 = weight_out_53[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_3 = weight_out_53[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_4 = weight_out_53[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_5 = weight_out_53[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_6 = weight_out_53[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_53_7 = weight_out_53[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_497 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_53_1 : read_data_53_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_498 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_53_2 : _GEN_497; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_499 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_53_3 : _GEN_498; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_500 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_53_4 : _GEN_499; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_501 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_53_5 : _GEN_500; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_502 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_53_6 : _GEN_501; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_53 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_53_7 : _GEN_502; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_54 = buf_unit_6_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_54_0 = weight_out_54[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_1 = weight_out_54[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_2 = weight_out_54[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_3 = weight_out_54[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_4 = weight_out_54[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_5 = weight_out_54[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_6 = weight_out_54[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_54_7 = weight_out_54[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_505 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_54_1 : read_data_54_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_506 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_54_2 : _GEN_505; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_507 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_54_3 : _GEN_506; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_508 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_54_4 : _GEN_507; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_509 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_54_5 : _GEN_508; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_510 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_54_6 : _GEN_509; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_54 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_54_7 : _GEN_510; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_55 = buf_unit_6_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_55_0 = weight_out_55[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_1 = weight_out_55[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_2 = weight_out_55[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_3 = weight_out_55[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_4 = weight_out_55[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_5 = weight_out_55[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_6 = weight_out_55[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_55_7 = weight_out_55[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_513 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_55_1 : read_data_55_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_514 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_55_2 : _GEN_513; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_515 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_55_3 : _GEN_514; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_516 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_55_4 : _GEN_515; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_517 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_55_5 : _GEN_516; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_518 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_55_6 : _GEN_517; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_55 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_55_7 : _GEN_518; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_56 = buf_unit_7_io_weight_out_0; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_56_0 = weight_out_56[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_1 = weight_out_56[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_2 = weight_out_56[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_3 = weight_out_56[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_4 = weight_out_56[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_5 = weight_out_56[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_6 = weight_out_56[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_56_7 = weight_out_56[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_521 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_56_1 : read_data_56_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_522 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_56_2 : _GEN_521; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_523 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_56_3 : _GEN_522; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_524 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_56_4 : _GEN_523; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_525 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_56_5 : _GEN_524; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_526 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_56_6 : _GEN_525; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_56 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_56_7 : _GEN_526; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_57 = buf_unit_7_io_weight_out_1; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_57_0 = weight_out_57[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_1 = weight_out_57[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_2 = weight_out_57[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_3 = weight_out_57[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_4 = weight_out_57[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_5 = weight_out_57[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_6 = weight_out_57[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_57_7 = weight_out_57[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_529 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_57_1 : read_data_57_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_530 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_57_2 : _GEN_529; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_531 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_57_3 : _GEN_530; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_532 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_57_4 : _GEN_531; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_533 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_57_5 : _GEN_532; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_534 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_57_6 : _GEN_533; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_57 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_57_7 : _GEN_534; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_58 = buf_unit_7_io_weight_out_2; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_58_0 = weight_out_58[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_1 = weight_out_58[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_2 = weight_out_58[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_3 = weight_out_58[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_4 = weight_out_58[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_5 = weight_out_58[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_6 = weight_out_58[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_58_7 = weight_out_58[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_537 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_58_1 : read_data_58_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_538 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_58_2 : _GEN_537; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_539 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_58_3 : _GEN_538; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_540 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_58_4 : _GEN_539; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_541 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_58_5 : _GEN_540; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_542 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_58_6 : _GEN_541; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_58 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_58_7 : _GEN_542; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_59 = buf_unit_7_io_weight_out_3; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_59_0 = weight_out_59[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_1 = weight_out_59[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_2 = weight_out_59[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_3 = weight_out_59[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_4 = weight_out_59[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_5 = weight_out_59[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_6 = weight_out_59[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_59_7 = weight_out_59[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_545 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_59_1 : read_data_59_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_546 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_59_2 : _GEN_545; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_547 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_59_3 : _GEN_546; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_548 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_59_4 : _GEN_547; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_549 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_59_5 : _GEN_548; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_550 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_59_6 : _GEN_549; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_59 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_59_7 : _GEN_550; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_60 = buf_unit_7_io_weight_out_4; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_60_0 = weight_out_60[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_1 = weight_out_60[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_2 = weight_out_60[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_3 = weight_out_60[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_4 = weight_out_60[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_5 = weight_out_60[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_6 = weight_out_60[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_60_7 = weight_out_60[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_553 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_60_1 : read_data_60_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_554 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_60_2 : _GEN_553; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_555 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_60_3 : _GEN_554; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_556 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_60_4 : _GEN_555; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_557 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_60_5 : _GEN_556; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_558 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_60_6 : _GEN_557; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_60 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_60_7 : _GEN_558; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_61 = buf_unit_7_io_weight_out_5; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_61_0 = weight_out_61[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_1 = weight_out_61[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_2 = weight_out_61[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_3 = weight_out_61[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_4 = weight_out_61[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_5 = weight_out_61[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_6 = weight_out_61[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_61_7 = weight_out_61[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_561 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_61_1 : read_data_61_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_562 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_61_2 : _GEN_561; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_563 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_61_3 : _GEN_562; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_564 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_61_4 : _GEN_563; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_565 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_61_5 : _GEN_564; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_566 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_61_6 : _GEN_565; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_61 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_61_7 : _GEN_566; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_62 = buf_unit_7_io_weight_out_6; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_62_0 = weight_out_62[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_1 = weight_out_62[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_2 = weight_out_62[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_3 = weight_out_62[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_4 = weight_out_62[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_5 = weight_out_62[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_6 = weight_out_62[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_62_7 = weight_out_62[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_569 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_62_1 : read_data_62_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_570 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_62_2 : _GEN_569; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_571 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_62_3 : _GEN_570; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_572 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_62_4 : _GEN_571; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_573 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_62_5 : _GEN_572; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_574 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_62_6 : _GEN_573; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_62 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_62_7 : _GEN_574; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] weight_out_63 = buf_unit_7_io_weight_out_7; // @[WeightBuffer.scala 66:24 81:38]
  wire [7:0] read_data_63_0 = weight_out_63[7:0]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_1 = weight_out_63[15:8]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_2 = weight_out_63[23:16]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_3 = weight_out_63[31:24]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_4 = weight_out_63[39:32]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_5 = weight_out_63[47:40]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_6 = weight_out_63[55:48]; // @[WeightBuffer.scala 71:43]
  wire [7:0] read_data_63_7 = weight_out_63[63:56]; // @[WeightBuffer.scala 71:43]
  wire [7:0] _GEN_577 = 3'h1 == io_sel_when_kernal_is_1 ? read_data_63_1 : read_data_63_0; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_578 = 3'h2 == io_sel_when_kernal_is_1 ? read_data_63_2 : _GEN_577; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_579 = 3'h3 == io_sel_when_kernal_is_1 ? read_data_63_3 : _GEN_578; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_580 = 3'h4 == io_sel_when_kernal_is_1 ? read_data_63_4 : _GEN_579; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_581 = 3'h5 == io_sel_when_kernal_is_1 ? read_data_63_5 : _GEN_580; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] _GEN_582 = 3'h6 == io_sel_when_kernal_is_1 ? read_data_63_6 : _GEN_581; // @[WeightBuffer.scala 73:{25,25}]
  wire [7:0] read_data_sel_63 = 3'h7 == io_sel_when_kernal_is_1 ? read_data_63_7 : _GEN_582; // @[WeightBuffer.scala 73:{25,25}]
  wire [71:0] _io_weight_out_0_T = {16'h0,read_data_sel_0,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_1_T = {16'h0,read_data_sel_1,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_2_T = {16'h0,read_data_sel_2,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_3_T = {16'h0,read_data_sel_3,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_4_T = {16'h0,read_data_sel_4,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_5_T = {16'h0,read_data_sel_5,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_6_T = {16'h0,read_data_sel_6,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_7_T = {16'h0,read_data_sel_7,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_8_T = {16'h0,read_data_sel_8,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_9_T = {16'h0,read_data_sel_9,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_10_T = {16'h0,read_data_sel_10,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_11_T = {16'h0,read_data_sel_11,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_12_T = {16'h0,read_data_sel_12,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_13_T = {16'h0,read_data_sel_13,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_14_T = {16'h0,read_data_sel_14,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_15_T = {16'h0,read_data_sel_15,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_16_T = {16'h0,read_data_sel_16,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_17_T = {16'h0,read_data_sel_17,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_18_T = {16'h0,read_data_sel_18,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_19_T = {16'h0,read_data_sel_19,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_20_T = {16'h0,read_data_sel_20,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_21_T = {16'h0,read_data_sel_21,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_22_T = {16'h0,read_data_sel_22,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_23_T = {16'h0,read_data_sel_23,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_24_T = {16'h0,read_data_sel_24,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_25_T = {16'h0,read_data_sel_25,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_26_T = {16'h0,read_data_sel_26,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_27_T = {16'h0,read_data_sel_27,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_28_T = {16'h0,read_data_sel_28,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_29_T = {16'h0,read_data_sel_29,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_30_T = {16'h0,read_data_sel_30,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_31_T = {16'h0,read_data_sel_31,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_32_T = {16'h0,read_data_sel_32,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_33_T = {16'h0,read_data_sel_33,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_34_T = {16'h0,read_data_sel_34,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_35_T = {16'h0,read_data_sel_35,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_36_T = {16'h0,read_data_sel_36,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_37_T = {16'h0,read_data_sel_37,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_38_T = {16'h0,read_data_sel_38,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_39_T = {16'h0,read_data_sel_39,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_40_T = {16'h0,read_data_sel_40,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_41_T = {16'h0,read_data_sel_41,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_42_T = {16'h0,read_data_sel_42,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_43_T = {16'h0,read_data_sel_43,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_44_T = {16'h0,read_data_sel_44,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_45_T = {16'h0,read_data_sel_45,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_46_T = {16'h0,read_data_sel_46,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_47_T = {16'h0,read_data_sel_47,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_48_T = {16'h0,read_data_sel_48,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_49_T = {16'h0,read_data_sel_49,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_50_T = {16'h0,read_data_sel_50,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_51_T = {16'h0,read_data_sel_51,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_52_T = {16'h0,read_data_sel_52,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_53_T = {16'h0,read_data_sel_53,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_54_T = {16'h0,read_data_sel_54,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_55_T = {16'h0,read_data_sel_55,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_56_T = {16'h0,read_data_sel_56,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_57_T = {16'h0,read_data_sel_57,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_58_T = {16'h0,read_data_sel_58,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_59_T = {16'h0,read_data_sel_59,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_60_T = {16'h0,read_data_sel_60,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_61_T = {16'h0,read_data_sel_61,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_62_T = {16'h0,read_data_sel_62,48'h0}; // @[Cat.scala 33:92]
  wire [71:0] _io_weight_out_63_T = {16'h0,read_data_sel_63,48'h0}; // @[Cat.scala 33:92]
  w_buffer_unit buf_unit_0 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_0_clock),
    .io_write_addr_0(buf_unit_0_io_write_addr_0),
    .io_write_addr_1(buf_unit_0_io_write_addr_1),
    .io_write_addr_2(buf_unit_0_io_write_addr_2),
    .io_write_addr_3(buf_unit_0_io_write_addr_3),
    .io_write_addr_4(buf_unit_0_io_write_addr_4),
    .io_write_addr_5(buf_unit_0_io_write_addr_5),
    .io_write_addr_6(buf_unit_0_io_write_addr_6),
    .io_write_addr_7(buf_unit_0_io_write_addr_7),
    .io_write_en_0(buf_unit_0_io_write_en_0),
    .io_write_en_1(buf_unit_0_io_write_en_1),
    .io_write_en_2(buf_unit_0_io_write_en_2),
    .io_write_en_3(buf_unit_0_io_write_en_3),
    .io_write_en_4(buf_unit_0_io_write_en_4),
    .io_write_en_5(buf_unit_0_io_write_en_5),
    .io_write_en_6(buf_unit_0_io_write_en_6),
    .io_write_en_7(buf_unit_0_io_write_en_7),
    .io_weight_in(buf_unit_0_io_weight_in),
    .io_read_addr(buf_unit_0_io_read_addr),
    .io_weight_out_0(buf_unit_0_io_weight_out_0),
    .io_weight_out_1(buf_unit_0_io_weight_out_1),
    .io_weight_out_2(buf_unit_0_io_weight_out_2),
    .io_weight_out_3(buf_unit_0_io_weight_out_3),
    .io_weight_out_4(buf_unit_0_io_weight_out_4),
    .io_weight_out_5(buf_unit_0_io_weight_out_5),
    .io_weight_out_6(buf_unit_0_io_weight_out_6),
    .io_weight_out_7(buf_unit_0_io_weight_out_7)
  );
  w_buffer_unit buf_unit_1 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_1_clock),
    .io_write_addr_0(buf_unit_1_io_write_addr_0),
    .io_write_addr_1(buf_unit_1_io_write_addr_1),
    .io_write_addr_2(buf_unit_1_io_write_addr_2),
    .io_write_addr_3(buf_unit_1_io_write_addr_3),
    .io_write_addr_4(buf_unit_1_io_write_addr_4),
    .io_write_addr_5(buf_unit_1_io_write_addr_5),
    .io_write_addr_6(buf_unit_1_io_write_addr_6),
    .io_write_addr_7(buf_unit_1_io_write_addr_7),
    .io_write_en_0(buf_unit_1_io_write_en_0),
    .io_write_en_1(buf_unit_1_io_write_en_1),
    .io_write_en_2(buf_unit_1_io_write_en_2),
    .io_write_en_3(buf_unit_1_io_write_en_3),
    .io_write_en_4(buf_unit_1_io_write_en_4),
    .io_write_en_5(buf_unit_1_io_write_en_5),
    .io_write_en_6(buf_unit_1_io_write_en_6),
    .io_write_en_7(buf_unit_1_io_write_en_7),
    .io_weight_in(buf_unit_1_io_weight_in),
    .io_read_addr(buf_unit_1_io_read_addr),
    .io_weight_out_0(buf_unit_1_io_weight_out_0),
    .io_weight_out_1(buf_unit_1_io_weight_out_1),
    .io_weight_out_2(buf_unit_1_io_weight_out_2),
    .io_weight_out_3(buf_unit_1_io_weight_out_3),
    .io_weight_out_4(buf_unit_1_io_weight_out_4),
    .io_weight_out_5(buf_unit_1_io_weight_out_5),
    .io_weight_out_6(buf_unit_1_io_weight_out_6),
    .io_weight_out_7(buf_unit_1_io_weight_out_7)
  );
  w_buffer_unit buf_unit_2 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_2_clock),
    .io_write_addr_0(buf_unit_2_io_write_addr_0),
    .io_write_addr_1(buf_unit_2_io_write_addr_1),
    .io_write_addr_2(buf_unit_2_io_write_addr_2),
    .io_write_addr_3(buf_unit_2_io_write_addr_3),
    .io_write_addr_4(buf_unit_2_io_write_addr_4),
    .io_write_addr_5(buf_unit_2_io_write_addr_5),
    .io_write_addr_6(buf_unit_2_io_write_addr_6),
    .io_write_addr_7(buf_unit_2_io_write_addr_7),
    .io_write_en_0(buf_unit_2_io_write_en_0),
    .io_write_en_1(buf_unit_2_io_write_en_1),
    .io_write_en_2(buf_unit_2_io_write_en_2),
    .io_write_en_3(buf_unit_2_io_write_en_3),
    .io_write_en_4(buf_unit_2_io_write_en_4),
    .io_write_en_5(buf_unit_2_io_write_en_5),
    .io_write_en_6(buf_unit_2_io_write_en_6),
    .io_write_en_7(buf_unit_2_io_write_en_7),
    .io_weight_in(buf_unit_2_io_weight_in),
    .io_read_addr(buf_unit_2_io_read_addr),
    .io_weight_out_0(buf_unit_2_io_weight_out_0),
    .io_weight_out_1(buf_unit_2_io_weight_out_1),
    .io_weight_out_2(buf_unit_2_io_weight_out_2),
    .io_weight_out_3(buf_unit_2_io_weight_out_3),
    .io_weight_out_4(buf_unit_2_io_weight_out_4),
    .io_weight_out_5(buf_unit_2_io_weight_out_5),
    .io_weight_out_6(buf_unit_2_io_weight_out_6),
    .io_weight_out_7(buf_unit_2_io_weight_out_7)
  );
  w_buffer_unit buf_unit_3 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_3_clock),
    .io_write_addr_0(buf_unit_3_io_write_addr_0),
    .io_write_addr_1(buf_unit_3_io_write_addr_1),
    .io_write_addr_2(buf_unit_3_io_write_addr_2),
    .io_write_addr_3(buf_unit_3_io_write_addr_3),
    .io_write_addr_4(buf_unit_3_io_write_addr_4),
    .io_write_addr_5(buf_unit_3_io_write_addr_5),
    .io_write_addr_6(buf_unit_3_io_write_addr_6),
    .io_write_addr_7(buf_unit_3_io_write_addr_7),
    .io_write_en_0(buf_unit_3_io_write_en_0),
    .io_write_en_1(buf_unit_3_io_write_en_1),
    .io_write_en_2(buf_unit_3_io_write_en_2),
    .io_write_en_3(buf_unit_3_io_write_en_3),
    .io_write_en_4(buf_unit_3_io_write_en_4),
    .io_write_en_5(buf_unit_3_io_write_en_5),
    .io_write_en_6(buf_unit_3_io_write_en_6),
    .io_write_en_7(buf_unit_3_io_write_en_7),
    .io_weight_in(buf_unit_3_io_weight_in),
    .io_read_addr(buf_unit_3_io_read_addr),
    .io_weight_out_0(buf_unit_3_io_weight_out_0),
    .io_weight_out_1(buf_unit_3_io_weight_out_1),
    .io_weight_out_2(buf_unit_3_io_weight_out_2),
    .io_weight_out_3(buf_unit_3_io_weight_out_3),
    .io_weight_out_4(buf_unit_3_io_weight_out_4),
    .io_weight_out_5(buf_unit_3_io_weight_out_5),
    .io_weight_out_6(buf_unit_3_io_weight_out_6),
    .io_weight_out_7(buf_unit_3_io_weight_out_7)
  );
  w_buffer_unit buf_unit_4 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_4_clock),
    .io_write_addr_0(buf_unit_4_io_write_addr_0),
    .io_write_addr_1(buf_unit_4_io_write_addr_1),
    .io_write_addr_2(buf_unit_4_io_write_addr_2),
    .io_write_addr_3(buf_unit_4_io_write_addr_3),
    .io_write_addr_4(buf_unit_4_io_write_addr_4),
    .io_write_addr_5(buf_unit_4_io_write_addr_5),
    .io_write_addr_6(buf_unit_4_io_write_addr_6),
    .io_write_addr_7(buf_unit_4_io_write_addr_7),
    .io_write_en_0(buf_unit_4_io_write_en_0),
    .io_write_en_1(buf_unit_4_io_write_en_1),
    .io_write_en_2(buf_unit_4_io_write_en_2),
    .io_write_en_3(buf_unit_4_io_write_en_3),
    .io_write_en_4(buf_unit_4_io_write_en_4),
    .io_write_en_5(buf_unit_4_io_write_en_5),
    .io_write_en_6(buf_unit_4_io_write_en_6),
    .io_write_en_7(buf_unit_4_io_write_en_7),
    .io_weight_in(buf_unit_4_io_weight_in),
    .io_read_addr(buf_unit_4_io_read_addr),
    .io_weight_out_0(buf_unit_4_io_weight_out_0),
    .io_weight_out_1(buf_unit_4_io_weight_out_1),
    .io_weight_out_2(buf_unit_4_io_weight_out_2),
    .io_weight_out_3(buf_unit_4_io_weight_out_3),
    .io_weight_out_4(buf_unit_4_io_weight_out_4),
    .io_weight_out_5(buf_unit_4_io_weight_out_5),
    .io_weight_out_6(buf_unit_4_io_weight_out_6),
    .io_weight_out_7(buf_unit_4_io_weight_out_7)
  );
  w_buffer_unit buf_unit_5 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_5_clock),
    .io_write_addr_0(buf_unit_5_io_write_addr_0),
    .io_write_addr_1(buf_unit_5_io_write_addr_1),
    .io_write_addr_2(buf_unit_5_io_write_addr_2),
    .io_write_addr_3(buf_unit_5_io_write_addr_3),
    .io_write_addr_4(buf_unit_5_io_write_addr_4),
    .io_write_addr_5(buf_unit_5_io_write_addr_5),
    .io_write_addr_6(buf_unit_5_io_write_addr_6),
    .io_write_addr_7(buf_unit_5_io_write_addr_7),
    .io_write_en_0(buf_unit_5_io_write_en_0),
    .io_write_en_1(buf_unit_5_io_write_en_1),
    .io_write_en_2(buf_unit_5_io_write_en_2),
    .io_write_en_3(buf_unit_5_io_write_en_3),
    .io_write_en_4(buf_unit_5_io_write_en_4),
    .io_write_en_5(buf_unit_5_io_write_en_5),
    .io_write_en_6(buf_unit_5_io_write_en_6),
    .io_write_en_7(buf_unit_5_io_write_en_7),
    .io_weight_in(buf_unit_5_io_weight_in),
    .io_read_addr(buf_unit_5_io_read_addr),
    .io_weight_out_0(buf_unit_5_io_weight_out_0),
    .io_weight_out_1(buf_unit_5_io_weight_out_1),
    .io_weight_out_2(buf_unit_5_io_weight_out_2),
    .io_weight_out_3(buf_unit_5_io_weight_out_3),
    .io_weight_out_4(buf_unit_5_io_weight_out_4),
    .io_weight_out_5(buf_unit_5_io_weight_out_5),
    .io_weight_out_6(buf_unit_5_io_weight_out_6),
    .io_weight_out_7(buf_unit_5_io_weight_out_7)
  );
  w_buffer_unit buf_unit_6 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_6_clock),
    .io_write_addr_0(buf_unit_6_io_write_addr_0),
    .io_write_addr_1(buf_unit_6_io_write_addr_1),
    .io_write_addr_2(buf_unit_6_io_write_addr_2),
    .io_write_addr_3(buf_unit_6_io_write_addr_3),
    .io_write_addr_4(buf_unit_6_io_write_addr_4),
    .io_write_addr_5(buf_unit_6_io_write_addr_5),
    .io_write_addr_6(buf_unit_6_io_write_addr_6),
    .io_write_addr_7(buf_unit_6_io_write_addr_7),
    .io_write_en_0(buf_unit_6_io_write_en_0),
    .io_write_en_1(buf_unit_6_io_write_en_1),
    .io_write_en_2(buf_unit_6_io_write_en_2),
    .io_write_en_3(buf_unit_6_io_write_en_3),
    .io_write_en_4(buf_unit_6_io_write_en_4),
    .io_write_en_5(buf_unit_6_io_write_en_5),
    .io_write_en_6(buf_unit_6_io_write_en_6),
    .io_write_en_7(buf_unit_6_io_write_en_7),
    .io_weight_in(buf_unit_6_io_weight_in),
    .io_read_addr(buf_unit_6_io_read_addr),
    .io_weight_out_0(buf_unit_6_io_weight_out_0),
    .io_weight_out_1(buf_unit_6_io_weight_out_1),
    .io_weight_out_2(buf_unit_6_io_weight_out_2),
    .io_weight_out_3(buf_unit_6_io_weight_out_3),
    .io_weight_out_4(buf_unit_6_io_weight_out_4),
    .io_weight_out_5(buf_unit_6_io_weight_out_5),
    .io_weight_out_6(buf_unit_6_io_weight_out_6),
    .io_weight_out_7(buf_unit_6_io_weight_out_7)
  );
  w_buffer_unit buf_unit_7 ( // @[WeightBuffer.scala 76:42]
    .clock(buf_unit_7_clock),
    .io_write_addr_0(buf_unit_7_io_write_addr_0),
    .io_write_addr_1(buf_unit_7_io_write_addr_1),
    .io_write_addr_2(buf_unit_7_io_write_addr_2),
    .io_write_addr_3(buf_unit_7_io_write_addr_3),
    .io_write_addr_4(buf_unit_7_io_write_addr_4),
    .io_write_addr_5(buf_unit_7_io_write_addr_5),
    .io_write_addr_6(buf_unit_7_io_write_addr_6),
    .io_write_addr_7(buf_unit_7_io_write_addr_7),
    .io_write_en_0(buf_unit_7_io_write_en_0),
    .io_write_en_1(buf_unit_7_io_write_en_1),
    .io_write_en_2(buf_unit_7_io_write_en_2),
    .io_write_en_3(buf_unit_7_io_write_en_3),
    .io_write_en_4(buf_unit_7_io_write_en_4),
    .io_write_en_5(buf_unit_7_io_write_en_5),
    .io_write_en_6(buf_unit_7_io_write_en_6),
    .io_write_en_7(buf_unit_7_io_write_en_7),
    .io_weight_in(buf_unit_7_io_weight_in),
    .io_read_addr(buf_unit_7_io_read_addr),
    .io_weight_out_0(buf_unit_7_io_weight_out_0),
    .io_weight_out_1(buf_unit_7_io_weight_out_1),
    .io_weight_out_2(buf_unit_7_io_weight_out_2),
    .io_weight_out_3(buf_unit_7_io_weight_out_3),
    .io_weight_out_4(buf_unit_7_io_weight_out_4),
    .io_weight_out_5(buf_unit_7_io_weight_out_5),
    .io_weight_out_6(buf_unit_7_io_weight_out_6),
    .io_weight_out_7(buf_unit_7_io_weight_out_7)
  );
  assign io_weight_out_0 = io_kernal ? weight_out_0 : _io_weight_out_0_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_1 = io_kernal ? weight_out_1 : _io_weight_out_1_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_2 = io_kernal ? weight_out_2 : _io_weight_out_2_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_3 = io_kernal ? weight_out_3 : _io_weight_out_3_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_4 = io_kernal ? weight_out_4 : _io_weight_out_4_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_5 = io_kernal ? weight_out_5 : _io_weight_out_5_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_6 = io_kernal ? weight_out_6 : _io_weight_out_6_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_7 = io_kernal ? weight_out_7 : _io_weight_out_7_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_8 = io_kernal ? weight_out_8 : _io_weight_out_8_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_9 = io_kernal ? weight_out_9 : _io_weight_out_9_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_10 = io_kernal ? weight_out_10 : _io_weight_out_10_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_11 = io_kernal ? weight_out_11 : _io_weight_out_11_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_12 = io_kernal ? weight_out_12 : _io_weight_out_12_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_13 = io_kernal ? weight_out_13 : _io_weight_out_13_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_14 = io_kernal ? weight_out_14 : _io_weight_out_14_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_15 = io_kernal ? weight_out_15 : _io_weight_out_15_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_16 = io_kernal ? weight_out_16 : _io_weight_out_16_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_17 = io_kernal ? weight_out_17 : _io_weight_out_17_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_18 = io_kernal ? weight_out_18 : _io_weight_out_18_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_19 = io_kernal ? weight_out_19 : _io_weight_out_19_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_20 = io_kernal ? weight_out_20 : _io_weight_out_20_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_21 = io_kernal ? weight_out_21 : _io_weight_out_21_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_22 = io_kernal ? weight_out_22 : _io_weight_out_22_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_23 = io_kernal ? weight_out_23 : _io_weight_out_23_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_24 = io_kernal ? weight_out_24 : _io_weight_out_24_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_25 = io_kernal ? weight_out_25 : _io_weight_out_25_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_26 = io_kernal ? weight_out_26 : _io_weight_out_26_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_27 = io_kernal ? weight_out_27 : _io_weight_out_27_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_28 = io_kernal ? weight_out_28 : _io_weight_out_28_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_29 = io_kernal ? weight_out_29 : _io_weight_out_29_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_30 = io_kernal ? weight_out_30 : _io_weight_out_30_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_31 = io_kernal ? weight_out_31 : _io_weight_out_31_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_32 = io_kernal ? weight_out_32 : _io_weight_out_32_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_33 = io_kernal ? weight_out_33 : _io_weight_out_33_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_34 = io_kernal ? weight_out_34 : _io_weight_out_34_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_35 = io_kernal ? weight_out_35 : _io_weight_out_35_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_36 = io_kernal ? weight_out_36 : _io_weight_out_36_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_37 = io_kernal ? weight_out_37 : _io_weight_out_37_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_38 = io_kernal ? weight_out_38 : _io_weight_out_38_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_39 = io_kernal ? weight_out_39 : _io_weight_out_39_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_40 = io_kernal ? weight_out_40 : _io_weight_out_40_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_41 = io_kernal ? weight_out_41 : _io_weight_out_41_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_42 = io_kernal ? weight_out_42 : _io_weight_out_42_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_43 = io_kernal ? weight_out_43 : _io_weight_out_43_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_44 = io_kernal ? weight_out_44 : _io_weight_out_44_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_45 = io_kernal ? weight_out_45 : _io_weight_out_45_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_46 = io_kernal ? weight_out_46 : _io_weight_out_46_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_47 = io_kernal ? weight_out_47 : _io_weight_out_47_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_48 = io_kernal ? weight_out_48 : _io_weight_out_48_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_49 = io_kernal ? weight_out_49 : _io_weight_out_49_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_50 = io_kernal ? weight_out_50 : _io_weight_out_50_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_51 = io_kernal ? weight_out_51 : _io_weight_out_51_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_52 = io_kernal ? weight_out_52 : _io_weight_out_52_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_53 = io_kernal ? weight_out_53 : _io_weight_out_53_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_54 = io_kernal ? weight_out_54 : _io_weight_out_54_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_55 = io_kernal ? weight_out_55 : _io_weight_out_55_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_56 = io_kernal ? weight_out_56 : _io_weight_out_56_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_57 = io_kernal ? weight_out_57 : _io_weight_out_57_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_58 = io_kernal ? weight_out_58 : _io_weight_out_58_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_59 = io_kernal ? weight_out_59 : _io_weight_out_59_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_60 = io_kernal ? weight_out_60 : _io_weight_out_60_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_61 = io_kernal ? weight_out_61 : _io_weight_out_61_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_62 = io_kernal ? weight_out_62 : _io_weight_out_62_T; // @[WeightBuffer.scala 82:45]
  assign io_weight_out_63 = io_kernal ? weight_out_63 : _io_weight_out_63_T; // @[WeightBuffer.scala 82:45]
  assign buf_unit_0_clock = clock;
  assign buf_unit_0_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_0_io_write_en_0 = ch_en_reg_0 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_1 = ch_en_reg_1 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_2 = ch_en_reg_2 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_3 = ch_en_reg_3 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_4 = ch_en_reg_4 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_5 = ch_en_reg_5 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_6 = ch_en_reg_6 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_write_en_7 = ch_en_reg_7 | force_write_0; // @[WeightBuffer.scala 80:56]
  assign buf_unit_0_io_weight_in = io_kernal ? w_data_when_k_is_3_0 : w_data_when_k_is_1_0; // @[WeightBuffer.scala 40:19]
  assign buf_unit_0_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_1_clock = clock;
  assign buf_unit_1_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_1_io_write_en_0 = ch_en_reg_0 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_1 = ch_en_reg_1 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_2 = ch_en_reg_2 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_3 = ch_en_reg_3 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_4 = ch_en_reg_4 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_5 = ch_en_reg_5 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_6 = ch_en_reg_6 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_write_en_7 = ch_en_reg_7 | force_write_1; // @[WeightBuffer.scala 80:56]
  assign buf_unit_1_io_weight_in = io_kernal ? w_data_when_k_is_3_1 : w_data_when_k_is_1_1; // @[WeightBuffer.scala 40:19]
  assign buf_unit_1_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_2_clock = clock;
  assign buf_unit_2_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_2_io_write_en_0 = ch_en_reg_0 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_1 = ch_en_reg_1 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_2 = ch_en_reg_2 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_3 = ch_en_reg_3 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_4 = ch_en_reg_4 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_5 = ch_en_reg_5 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_6 = ch_en_reg_6 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_write_en_7 = ch_en_reg_7 | force_write_2; // @[WeightBuffer.scala 80:56]
  assign buf_unit_2_io_weight_in = io_kernal ? w_data_when_k_is_3_2 : w_data_when_k_is_1_2; // @[WeightBuffer.scala 40:19]
  assign buf_unit_2_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_3_clock = clock;
  assign buf_unit_3_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_3_io_write_en_0 = ch_en_reg_0 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_1 = ch_en_reg_1 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_2 = ch_en_reg_2 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_3 = ch_en_reg_3 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_4 = ch_en_reg_4 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_5 = ch_en_reg_5 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_6 = ch_en_reg_6 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_write_en_7 = ch_en_reg_7 | force_write_3; // @[WeightBuffer.scala 80:56]
  assign buf_unit_3_io_weight_in = io_kernal ? w_data_when_k_is_3_3 : w_data_when_k_is_1_3; // @[WeightBuffer.scala 40:19]
  assign buf_unit_3_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_4_clock = clock;
  assign buf_unit_4_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_4_io_write_en_0 = ch_en_reg_0 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_1 = ch_en_reg_1 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_2 = ch_en_reg_2 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_3 = ch_en_reg_3 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_4 = ch_en_reg_4 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_5 = ch_en_reg_5 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_6 = ch_en_reg_6 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_write_en_7 = ch_en_reg_7 | force_write_4; // @[WeightBuffer.scala 80:56]
  assign buf_unit_4_io_weight_in = io_kernal ? w_data_when_k_is_3_4 : w_data_when_k_is_1_4; // @[WeightBuffer.scala 40:19]
  assign buf_unit_4_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_5_clock = clock;
  assign buf_unit_5_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_5_io_write_en_0 = ch_en_reg_0 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_1 = ch_en_reg_1 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_2 = ch_en_reg_2 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_3 = ch_en_reg_3 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_4 = ch_en_reg_4 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_5 = ch_en_reg_5 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_6 = ch_en_reg_6 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_write_en_7 = ch_en_reg_7 | force_write_5; // @[WeightBuffer.scala 80:56]
  assign buf_unit_5_io_weight_in = io_kernal ? w_data_when_k_is_3_5 : w_data_when_k_is_1_5; // @[WeightBuffer.scala 40:19]
  assign buf_unit_5_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_6_clock = clock;
  assign buf_unit_6_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_6_io_write_en_0 = ch_en_reg_0 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_1 = ch_en_reg_1 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_2 = ch_en_reg_2 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_3 = ch_en_reg_3 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_4 = ch_en_reg_4 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_5 = ch_en_reg_5 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_6 = ch_en_reg_6 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_write_en_7 = ch_en_reg_7 | force_write_6; // @[WeightBuffer.scala 80:56]
  assign buf_unit_6_io_weight_in = io_kernal ? w_data_when_k_is_3_6 : w_data_when_k_is_1_6; // @[WeightBuffer.scala 40:19]
  assign buf_unit_6_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  assign buf_unit_7_clock = clock;
  assign buf_unit_7_io_write_addr_0 = ch_cnt_0; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_1 = ch_cnt_1; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_2 = ch_cnt_2; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_3 = ch_cnt_3; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_4 = ch_cnt_4; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_5 = ch_cnt_5; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_6 = ch_cnt_6; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_addr_7 = ch_cnt_7; // @[WeightBuffer.scala 79:42]
  assign buf_unit_7_io_write_en_0 = ch_en_reg_0 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_1 = ch_en_reg_1 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_2 = ch_en_reg_2 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_3 = ch_en_reg_3 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_4 = ch_en_reg_4 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_5 = ch_en_reg_5 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_6 = ch_en_reg_6 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_write_en_7 = ch_en_reg_7 | force_write_7; // @[WeightBuffer.scala 80:56]
  assign buf_unit_7_io_weight_in = io_kernal ? w_data_when_k_is_3_7 : w_data_when_k_is_1_7; // @[WeightBuffer.scala 40:19]
  assign buf_unit_7_io_read_addr = io_read_addr; // @[WeightBuffer.scala 85:34]
  always @(posedge clock) begin
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_0 <= io_in_0; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_1 <= temp_0_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_2 <= temp_0_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_3 <= temp_0_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_4 <= temp_0_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_5 <= temp_0_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_6 <= temp_0_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_7 <= temp_0_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_0_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_0_8 <= temp_0_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_0 <= io_in_1; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_1 <= temp_1_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_2 <= temp_1_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_3 <= temp_1_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_4 <= temp_1_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_5 <= temp_1_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_6 <= temp_1_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_7 <= temp_1_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_1_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_1_8 <= temp_1_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_0 <= io_in_2; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_1 <= temp_2_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_2 <= temp_2_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_3 <= temp_2_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_4 <= temp_2_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_5 <= temp_2_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_6 <= temp_2_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_7 <= temp_2_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_2_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_2_8 <= temp_2_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_0 <= io_in_3; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_1 <= temp_3_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_2 <= temp_3_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_3 <= temp_3_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_4 <= temp_3_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_5 <= temp_3_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_6 <= temp_3_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_7 <= temp_3_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_3_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_3_8 <= temp_3_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_0 <= io_in_4; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_1 <= temp_4_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_2 <= temp_4_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_3 <= temp_4_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_4 <= temp_4_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_5 <= temp_4_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_6 <= temp_4_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_7 <= temp_4_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_4_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_4_8 <= temp_4_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_0 <= io_in_5; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_1 <= temp_5_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_2 <= temp_5_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_3 <= temp_5_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_4 <= temp_5_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_5 <= temp_5_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_6 <= temp_5_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_7 <= temp_5_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_5_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_5_8 <= temp_5_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_0 <= io_in_6; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_1 <= temp_6_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_2 <= temp_6_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_3 <= temp_6_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_4 <= temp_6_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_5 <= temp_6_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_6 <= temp_6_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_7 <= temp_6_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_6_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_6_8 <= temp_6_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_0 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_0 <= io_in_7; // @[WeightBuffer.scala 23:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_1 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_1 <= temp_7_0; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_2 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_2 <= temp_7_1; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_3 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_3 <= temp_7_2; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_4 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_4 <= temp_7_3; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_5 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_5 <= temp_7_4; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_6 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_6 <= temp_7_5; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_7 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_7 <= temp_7_6; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 17:51]
      temp_7_8 <= 8'h0; // @[WeightBuffer.scala 17:51]
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 19:5]
      temp_7_8 <= temp_7_7; // @[WeightBuffer.scala 26:32]
    end
    if (reset) begin // @[WeightBuffer.scala 42:23]
      cnt9 <= 4'h0; // @[WeightBuffer.scala 42:23]
    end else if (rst) begin // @[WeightBuffer.scala 46:16]
      cnt9 <= 4'h0;
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 46:30]
      if (cnt9 == cnt9_max) begin // @[WeightBuffer.scala 46:52]
        cnt9 <= 4'h0;
      end else begin
        cnt9 <= _cnt9_T_2;
      end
    end
    if (reset) begin // @[WeightBuffer.scala 44:23]
      cnt8 <= 3'h0; // @[WeightBuffer.scala 44:23]
    end else if (rst) begin // @[WeightBuffer.scala 47:16]
      cnt8 <= 3'h0;
    end else if (io_bram_write_en) begin // @[WeightBuffer.scala 47:30]
      if (_cnt9_T) begin // @[WeightBuffer.scala 47:52]
        cnt8 <= _cnt8_T_4;
      end
    end
    ch_en_reg_0 <= io_bram_write_en & cnt8 == 3'h0 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_1 <= io_bram_write_en & cnt8 == 3'h1 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_2 <= io_bram_write_en & cnt8 == 3'h2 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_3 <= io_bram_write_en & cnt8 == 3'h3 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_4 <= io_bram_write_en & cnt8 == 3'h4 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_5 <= io_bram_write_en & cnt8 == 3'h5 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_6 <= io_bram_write_en & cnt8 == 3'h6 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    ch_en_reg_7 <= io_bram_write_en & _cnt8_T_1 & _cnt9_T; // @[WeightBuffer.scala 51:56]
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_0 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_0 <= 7'h0;
    end else if (ch_en_reg_0) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_0 <= _ch_cnt_0_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_1 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_1 <= 7'h0;
    end else if (ch_en_reg_1) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_1 <= _ch_cnt_1_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_2 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_2 <= 7'h0;
    end else if (ch_en_reg_2) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_2 <= _ch_cnt_2_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_3 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_3 <= 7'h0;
    end else if (ch_en_reg_3) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_3 <= _ch_cnt_3_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_4 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_4 <= 7'h0;
    end else if (ch_en_reg_4) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_4 <= _ch_cnt_4_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_5 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_5 <= 7'h0;
    end else if (ch_en_reg_5) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_5 <= _ch_cnt_5_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_6 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_6 <= 7'h0;
    end else if (ch_en_reg_6) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_6 <= _ch_cnt_6_T_1;
    end
    if (reset) begin // @[WeightBuffer.scala 55:40]
      ch_cnt_7 <= 7'h0; // @[WeightBuffer.scala 55:40]
    end else if (rst) begin // @[WeightBuffer.scala 57:25]
      ch_cnt_7 <= 7'h0;
    end else if (ch_en_reg_7) begin // @[WeightBuffer.scala 57:39]
      ch_cnt_7 <= _ch_cnt_7_T_1;
    end
    if (reset) begin // @[utils.scala 19:16]
      bram_write_en_downedge_REG <= 1'h0; // @[utils.scala 19:16]
    end else begin
      bram_write_en_downedge_REG <= io_bram_write_en; // @[utils.scala 19:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  temp_0_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  temp_0_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  temp_0_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  temp_0_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  temp_0_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  temp_0_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  temp_0_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  temp_0_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  temp_1_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  temp_1_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  temp_1_2 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  temp_1_3 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  temp_1_4 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  temp_1_5 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  temp_1_6 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  temp_1_7 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  temp_1_8 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  temp_2_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  temp_2_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  temp_2_2 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  temp_2_3 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  temp_2_4 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  temp_2_5 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  temp_2_6 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  temp_2_7 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  temp_2_8 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  temp_3_0 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  temp_3_1 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  temp_3_2 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  temp_3_3 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  temp_3_4 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  temp_3_5 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  temp_3_6 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  temp_3_7 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  temp_3_8 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  temp_4_0 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  temp_4_1 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  temp_4_2 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  temp_4_3 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  temp_4_4 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  temp_4_5 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  temp_4_6 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  temp_4_7 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  temp_4_8 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  temp_5_0 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  temp_5_1 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  temp_5_2 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  temp_5_3 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  temp_5_4 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  temp_5_5 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  temp_5_6 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  temp_5_7 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  temp_5_8 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  temp_6_0 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  temp_6_1 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  temp_6_2 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  temp_6_3 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  temp_6_4 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  temp_6_5 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  temp_6_6 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  temp_6_7 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  temp_6_8 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  temp_7_0 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  temp_7_1 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  temp_7_2 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  temp_7_3 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  temp_7_4 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  temp_7_5 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  temp_7_6 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  temp_7_7 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  temp_7_8 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  cnt9 = _RAND_72[3:0];
  _RAND_73 = {1{`RANDOM}};
  cnt8 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  ch_en_reg_0 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  ch_en_reg_1 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  ch_en_reg_2 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  ch_en_reg_3 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  ch_en_reg_4 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  ch_en_reg_5 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  ch_en_reg_6 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  ch_en_reg_7 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  ch_cnt_0 = _RAND_82[6:0];
  _RAND_83 = {1{`RANDOM}};
  ch_cnt_1 = _RAND_83[6:0];
  _RAND_84 = {1{`RANDOM}};
  ch_cnt_2 = _RAND_84[6:0];
  _RAND_85 = {1{`RANDOM}};
  ch_cnt_3 = _RAND_85[6:0];
  _RAND_86 = {1{`RANDOM}};
  ch_cnt_4 = _RAND_86[6:0];
  _RAND_87 = {1{`RANDOM}};
  ch_cnt_5 = _RAND_87[6:0];
  _RAND_88 = {1{`RANDOM}};
  ch_cnt_6 = _RAND_88[6:0];
  _RAND_89 = {1{`RANDOM}};
  ch_cnt_7 = _RAND_89[6:0];
  _RAND_90 = {1{`RANDOM}};
  bram_write_en_downedge_REG = _RAND_90[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TPRAM_WRAP_80(
  input         clock,
  input         io_wen,
  input  [6:0]  io_waddr,
  input  [6:0]  io_raddr,
  input  [17:0] io_wdata,
  output [17:0] io_rdata
);
  wire  tpram_CLKA; // @[utils.scala 218:23]
  wire  tpram_CLKB; // @[utils.scala 218:23]
  wire  tpram_CENB; // @[utils.scala 218:23]
  wire  tpram_CENA; // @[utils.scala 218:23]
  wire [6:0] tpram_AB; // @[utils.scala 218:23]
  wire [6:0] tpram_AA; // @[utils.scala 218:23]
  wire [17:0] tpram_DB; // @[utils.scala 218:23]
  wire [17:0] tpram_QA; // @[utils.scala 218:23]
  TPRAM #(.DATA_WIDTH(18), .DEPTH(128), .RAM_STYLE_VAL("distributed")) tpram ( // @[utils.scala 218:23]
    .CLKA(tpram_CLKA),
    .CLKB(tpram_CLKB),
    .CENB(tpram_CENB),
    .CENA(tpram_CENA),
    .AB(tpram_AB),
    .AA(tpram_AA),
    .DB(tpram_DB),
    .QA(tpram_QA)
  );
  assign io_rdata = tpram_QA; // @[utils.scala 230:12]
  assign tpram_CLKA = clock; // @[utils.scala 222:19]
  assign tpram_CLKB = clock; // @[utils.scala 223:19]
  assign tpram_CENB = ~io_wen; // @[utils.scala 224:22]
  assign tpram_CENA = 1'h0; // @[utils.scala 225:22]
  assign tpram_AB = io_waddr; // @[utils.scala 226:17]
  assign tpram_AA = io_raddr; // @[utils.scala 227:17]
  assign tpram_DB = io_wdata; // @[utils.scala 228:17]
endmodule
module BiasBuffer(
  input         clock,
  input         reset,
  input         io_clear,
  input  [17:0] io_bias_in,
  input  [6:0]  io_bram_addr_read,
  input         io_bram_en_write,
  output [17:0] io_bias_data_0,
  output [17:0] io_bias_data_1,
  output [17:0] io_bias_data_2,
  output [17:0] io_bias_data_3,
  output [17:0] io_bias_data_4,
  output [17:0] io_bias_data_5,
  output [17:0] io_bias_data_6,
  output [17:0] io_bias_data_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  TPRAM_WRAP_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_1_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_1_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_1_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_1_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_1_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_2_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_2_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_2_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_2_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_2_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_3_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_3_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_3_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_3_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_3_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_4_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_4_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_4_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_4_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_4_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_5_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_5_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_5_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_5_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_5_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_6_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_6_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_6_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_6_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_6_io_rdata; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_7_io_wen; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_7_io_waddr; // @[utils.scala 237:100]
  wire [6:0] TPRAM_WRAP_7_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_7_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_7_io_rdata; // @[utils.scala 237:100]
  reg [2:0] cnt_8; // @[BiasBuffer.scala 14:24]
  reg [6:0] ch_cnt_0; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_1; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_2; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_3; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_4; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_5; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_6; // @[BiasBuffer.scala 15:21]
  reg [6:0] ch_cnt_7; // @[BiasBuffer.scala 15:21]
  reg  ch_en_reg_0; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_1; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_2; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_3; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_4; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_5; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_6; // @[BiasBuffer.scala 17:24]
  reg  ch_en_reg_7; // @[BiasBuffer.scala 17:24]
  wire  rst = io_clear | reset; // @[BiasBuffer.scala 18:24]
  wire [6:0] _ch_cnt_0_T_1 = ch_cnt_0 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_1_T_1 = ch_cnt_1 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_2_T_1 = ch_cnt_2 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_3_T_1 = ch_cnt_3 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_4_T_1 = ch_cnt_4 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_5_T_1 = ch_cnt_5 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_6_T_1 = ch_cnt_6 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [6:0] _ch_cnt_7_T_1 = ch_cnt_7 + 7'h1; // @[BiasBuffer.scala 22:64]
  wire [2:0] _cnt_8_T_1 = cnt_8 + 3'h1; // @[BiasBuffer.scala 24:56]
  TPRAM_WRAP_80 TPRAM_WRAP ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_clock),
    .io_wen(TPRAM_WRAP_io_wen),
    .io_waddr(TPRAM_WRAP_io_waddr),
    .io_raddr(TPRAM_WRAP_io_raddr),
    .io_wdata(TPRAM_WRAP_io_wdata),
    .io_rdata(TPRAM_WRAP_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_1 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_1_clock),
    .io_wen(TPRAM_WRAP_1_io_wen),
    .io_waddr(TPRAM_WRAP_1_io_waddr),
    .io_raddr(TPRAM_WRAP_1_io_raddr),
    .io_wdata(TPRAM_WRAP_1_io_wdata),
    .io_rdata(TPRAM_WRAP_1_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_2 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_2_clock),
    .io_wen(TPRAM_WRAP_2_io_wen),
    .io_waddr(TPRAM_WRAP_2_io_waddr),
    .io_raddr(TPRAM_WRAP_2_io_raddr),
    .io_wdata(TPRAM_WRAP_2_io_wdata),
    .io_rdata(TPRAM_WRAP_2_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_3 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_3_clock),
    .io_wen(TPRAM_WRAP_3_io_wen),
    .io_waddr(TPRAM_WRAP_3_io_waddr),
    .io_raddr(TPRAM_WRAP_3_io_raddr),
    .io_wdata(TPRAM_WRAP_3_io_wdata),
    .io_rdata(TPRAM_WRAP_3_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_4 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_4_clock),
    .io_wen(TPRAM_WRAP_4_io_wen),
    .io_waddr(TPRAM_WRAP_4_io_waddr),
    .io_raddr(TPRAM_WRAP_4_io_raddr),
    .io_wdata(TPRAM_WRAP_4_io_wdata),
    .io_rdata(TPRAM_WRAP_4_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_5 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_5_clock),
    .io_wen(TPRAM_WRAP_5_io_wen),
    .io_waddr(TPRAM_WRAP_5_io_waddr),
    .io_raddr(TPRAM_WRAP_5_io_raddr),
    .io_wdata(TPRAM_WRAP_5_io_wdata),
    .io_rdata(TPRAM_WRAP_5_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_6 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_6_clock),
    .io_wen(TPRAM_WRAP_6_io_wen),
    .io_waddr(TPRAM_WRAP_6_io_waddr),
    .io_raddr(TPRAM_WRAP_6_io_raddr),
    .io_wdata(TPRAM_WRAP_6_io_wdata),
    .io_rdata(TPRAM_WRAP_6_io_rdata)
  );
  TPRAM_WRAP_80 TPRAM_WRAP_7 ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_7_clock),
    .io_wen(TPRAM_WRAP_7_io_wen),
    .io_waddr(TPRAM_WRAP_7_io_waddr),
    .io_raddr(TPRAM_WRAP_7_io_raddr),
    .io_wdata(TPRAM_WRAP_7_io_wdata),
    .io_rdata(TPRAM_WRAP_7_io_rdata)
  );
  assign io_bias_data_0 = TPRAM_WRAP_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_1 = TPRAM_WRAP_1_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_2 = TPRAM_WRAP_2_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_3 = TPRAM_WRAP_3_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_4 = TPRAM_WRAP_4_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_5 = TPRAM_WRAP_5_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_6 = TPRAM_WRAP_6_io_rdata; // @[BiasBuffer.scala 34:25]
  assign io_bias_data_7 = TPRAM_WRAP_7_io_rdata; // @[BiasBuffer.scala 34:25]
  assign TPRAM_WRAP_clock = clock;
  assign TPRAM_WRAP_io_wen = io_bram_en_write & cnt_8 == 3'h0; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_io_waddr = ch_cnt_0; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_1_clock = clock;
  assign TPRAM_WRAP_1_io_wen = io_bram_en_write & cnt_8 == 3'h1; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_1_io_waddr = ch_cnt_1; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_1_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_1_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_2_clock = clock;
  assign TPRAM_WRAP_2_io_wen = io_bram_en_write & cnt_8 == 3'h2; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_2_io_waddr = ch_cnt_2; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_2_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_2_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_3_clock = clock;
  assign TPRAM_WRAP_3_io_wen = io_bram_en_write & cnt_8 == 3'h3; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_3_io_waddr = ch_cnt_3; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_3_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_3_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_4_clock = clock;
  assign TPRAM_WRAP_4_io_wen = io_bram_en_write & cnt_8 == 3'h4; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_4_io_waddr = ch_cnt_4; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_4_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_4_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_5_clock = clock;
  assign TPRAM_WRAP_5_io_wen = io_bram_en_write & cnt_8 == 3'h5; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_5_io_waddr = ch_cnt_5; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_5_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_5_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_6_clock = clock;
  assign TPRAM_WRAP_6_io_wen = io_bram_en_write & cnt_8 == 3'h6; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_6_io_waddr = ch_cnt_6; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_6_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_6_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  assign TPRAM_WRAP_7_clock = clock;
  assign TPRAM_WRAP_7_io_wen = io_bram_en_write & cnt_8 == 3'h7; // @[BiasBuffer.scala 20:38]
  assign TPRAM_WRAP_7_io_waddr = ch_cnt_7; // @[BiasBuffer.scala 31:22]
  assign TPRAM_WRAP_7_io_raddr = io_bram_addr_read; // @[BiasBuffer.scala 32:22]
  assign TPRAM_WRAP_7_io_wdata = io_bias_in; // @[BiasBuffer.scala 33:22]
  always @(posedge clock) begin
    if (reset) begin // @[BiasBuffer.scala 14:24]
      cnt_8 <= 3'h0; // @[BiasBuffer.scala 14:24]
    end else if (rst) begin // @[BiasBuffer.scala 24:17]
      cnt_8 <= 3'h0;
    end else if (io_bram_en_write) begin // @[BiasBuffer.scala 24:31]
      cnt_8 <= _cnt_8_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_0 <= 7'h0;
    end else if (ch_en_reg_0) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_0 <= _ch_cnt_0_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_1 <= 7'h0;
    end else if (ch_en_reg_1) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_1 <= _ch_cnt_1_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_2 <= 7'h0;
    end else if (ch_en_reg_2) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_2 <= _ch_cnt_2_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_3 <= 7'h0;
    end else if (ch_en_reg_3) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_3 <= _ch_cnt_3_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_4 <= 7'h0;
    end else if (ch_en_reg_4) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_4 <= _ch_cnt_4_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_5 <= 7'h0;
    end else if (ch_en_reg_5) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_5 <= _ch_cnt_5_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_6 <= 7'h0;
    end else if (ch_en_reg_6) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_6 <= _ch_cnt_6_T_1;
    end
    if (rst) begin // @[BiasBuffer.scala 22:25]
      ch_cnt_7 <= 7'h0;
    end else if (ch_en_reg_7) begin // @[BiasBuffer.scala 22:39]
      ch_cnt_7 <= _ch_cnt_7_T_1;
    end
    ch_en_reg_0 <= io_bram_en_write & cnt_8 == 3'h0; // @[BiasBuffer.scala 20:38]
    ch_en_reg_1 <= io_bram_en_write & cnt_8 == 3'h1; // @[BiasBuffer.scala 20:38]
    ch_en_reg_2 <= io_bram_en_write & cnt_8 == 3'h2; // @[BiasBuffer.scala 20:38]
    ch_en_reg_3 <= io_bram_en_write & cnt_8 == 3'h3; // @[BiasBuffer.scala 20:38]
    ch_en_reg_4 <= io_bram_en_write & cnt_8 == 3'h4; // @[BiasBuffer.scala 20:38]
    ch_en_reg_5 <= io_bram_en_write & cnt_8 == 3'h5; // @[BiasBuffer.scala 20:38]
    ch_en_reg_6 <= io_bram_en_write & cnt_8 == 3'h6; // @[BiasBuffer.scala 20:38]
    ch_en_reg_7 <= io_bram_en_write & cnt_8 == 3'h7; // @[BiasBuffer.scala 20:38]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt_8 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  ch_cnt_0 = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  ch_cnt_1 = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  ch_cnt_2 = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  ch_cnt_3 = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  ch_cnt_4 = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  ch_cnt_5 = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  ch_cnt_6 = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  ch_cnt_7 = _RAND_8[6:0];
  _RAND_9 = {1{`RANDOM}};
  ch_en_reg_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ch_en_reg_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ch_en_reg_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ch_en_reg_3 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ch_en_reg_4 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ch_en_reg_5 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ch_en_reg_6 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ch_en_reg_7 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cal_sub_zero_point(
  input        clock,
  input        reset,
  input  [7:0] io_zero_point,
  input  [7:0] io_data_in,
  output [7:0] io_data_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] out; // @[quant.scala 94:22]
  wire [7:0] _out_T_2 = $signed(io_data_in) - $signed(io_zero_point); // @[quant.scala 95:15]
  assign io_data_out = out; // @[quant.scala 96:24]
  always @(posedge clock) begin
    if (reset) begin // @[quant.scala 94:22]
      out <= 8'sh0; // @[quant.scala 94:22]
    end else begin
      out <= _out_T_2; // @[quant.scala 95:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module sub_zero_point(
  input        clock,
  input        reset,
  input  [7:0] io_zero_point,
  input  [7:0] io_data_in_0,
  input  [7:0] io_data_in_1,
  input  [7:0] io_data_in_2,
  input  [7:0] io_data_in_3,
  input  [7:0] io_data_in_4,
  input  [7:0] io_data_in_5,
  input  [7:0] io_data_in_6,
  input  [7:0] io_data_in_7,
  input  [7:0] io_data_in_8,
  input  [7:0] io_data_in_9,
  input  [7:0] io_data_in_10,
  input  [7:0] io_data_in_11,
  input  [7:0] io_data_in_12,
  input  [7:0] io_data_in_13,
  input  [7:0] io_data_in_14,
  input  [7:0] io_data_in_15,
  input  [7:0] io_data_in_16,
  input  [7:0] io_data_in_17,
  input  [7:0] io_data_in_18,
  input  [7:0] io_data_in_19,
  input  [7:0] io_data_in_20,
  input  [7:0] io_data_in_21,
  input  [7:0] io_data_in_22,
  input  [7:0] io_data_in_23,
  input  [7:0] io_data_in_24,
  input  [7:0] io_data_in_25,
  input  [7:0] io_data_in_26,
  input  [7:0] io_data_in_27,
  input  [7:0] io_data_in_28,
  input  [7:0] io_data_in_29,
  input  [7:0] io_data_in_30,
  input  [7:0] io_data_in_31,
  output [7:0] io_data_out_0,
  output [7:0] io_data_out_1,
  output [7:0] io_data_out_2,
  output [7:0] io_data_out_3,
  output [7:0] io_data_out_4,
  output [7:0] io_data_out_5,
  output [7:0] io_data_out_6,
  output [7:0] io_data_out_7,
  output [7:0] io_data_out_8,
  output [7:0] io_data_out_9,
  output [7:0] io_data_out_10,
  output [7:0] io_data_out_11,
  output [7:0] io_data_out_12,
  output [7:0] io_data_out_13,
  output [7:0] io_data_out_14,
  output [7:0] io_data_out_15,
  output [7:0] io_data_out_16,
  output [7:0] io_data_out_17,
  output [7:0] io_data_out_18,
  output [7:0] io_data_out_19,
  output [7:0] io_data_out_20,
  output [7:0] io_data_out_21,
  output [7:0] io_data_out_22,
  output [7:0] io_data_out_23,
  output [7:0] io_data_out_24,
  output [7:0] io_data_out_25,
  output [7:0] io_data_out_26,
  output [7:0] io_data_out_27,
  output [7:0] io_data_out_28,
  output [7:0] io_data_out_29,
  output [7:0] io_data_out_30,
  output [7:0] io_data_out_31
);
  wire  unit_0_clock; // @[quant.scala 78:52]
  wire  unit_0_reset; // @[quant.scala 78:52]
  wire [7:0] unit_0_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_0_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_0_io_data_out; // @[quant.scala 78:52]
  wire  unit_1_clock; // @[quant.scala 78:52]
  wire  unit_1_reset; // @[quant.scala 78:52]
  wire [7:0] unit_1_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_1_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_1_io_data_out; // @[quant.scala 78:52]
  wire  unit_2_clock; // @[quant.scala 78:52]
  wire  unit_2_reset; // @[quant.scala 78:52]
  wire [7:0] unit_2_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_2_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_2_io_data_out; // @[quant.scala 78:52]
  wire  unit_3_clock; // @[quant.scala 78:52]
  wire  unit_3_reset; // @[quant.scala 78:52]
  wire [7:0] unit_3_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_3_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_3_io_data_out; // @[quant.scala 78:52]
  wire  unit_4_clock; // @[quant.scala 78:52]
  wire  unit_4_reset; // @[quant.scala 78:52]
  wire [7:0] unit_4_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_4_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_4_io_data_out; // @[quant.scala 78:52]
  wire  unit_5_clock; // @[quant.scala 78:52]
  wire  unit_5_reset; // @[quant.scala 78:52]
  wire [7:0] unit_5_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_5_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_5_io_data_out; // @[quant.scala 78:52]
  wire  unit_6_clock; // @[quant.scala 78:52]
  wire  unit_6_reset; // @[quant.scala 78:52]
  wire [7:0] unit_6_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_6_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_6_io_data_out; // @[quant.scala 78:52]
  wire  unit_7_clock; // @[quant.scala 78:52]
  wire  unit_7_reset; // @[quant.scala 78:52]
  wire [7:0] unit_7_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_7_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_7_io_data_out; // @[quant.scala 78:52]
  wire  unit_8_clock; // @[quant.scala 78:52]
  wire  unit_8_reset; // @[quant.scala 78:52]
  wire [7:0] unit_8_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_8_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_8_io_data_out; // @[quant.scala 78:52]
  wire  unit_9_clock; // @[quant.scala 78:52]
  wire  unit_9_reset; // @[quant.scala 78:52]
  wire [7:0] unit_9_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_9_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_9_io_data_out; // @[quant.scala 78:52]
  wire  unit_10_clock; // @[quant.scala 78:52]
  wire  unit_10_reset; // @[quant.scala 78:52]
  wire [7:0] unit_10_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_10_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_10_io_data_out; // @[quant.scala 78:52]
  wire  unit_11_clock; // @[quant.scala 78:52]
  wire  unit_11_reset; // @[quant.scala 78:52]
  wire [7:0] unit_11_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_11_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_11_io_data_out; // @[quant.scala 78:52]
  wire  unit_12_clock; // @[quant.scala 78:52]
  wire  unit_12_reset; // @[quant.scala 78:52]
  wire [7:0] unit_12_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_12_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_12_io_data_out; // @[quant.scala 78:52]
  wire  unit_13_clock; // @[quant.scala 78:52]
  wire  unit_13_reset; // @[quant.scala 78:52]
  wire [7:0] unit_13_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_13_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_13_io_data_out; // @[quant.scala 78:52]
  wire  unit_14_clock; // @[quant.scala 78:52]
  wire  unit_14_reset; // @[quant.scala 78:52]
  wire [7:0] unit_14_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_14_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_14_io_data_out; // @[quant.scala 78:52]
  wire  unit_15_clock; // @[quant.scala 78:52]
  wire  unit_15_reset; // @[quant.scala 78:52]
  wire [7:0] unit_15_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_15_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_15_io_data_out; // @[quant.scala 78:52]
  wire  unit_16_clock; // @[quant.scala 78:52]
  wire  unit_16_reset; // @[quant.scala 78:52]
  wire [7:0] unit_16_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_16_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_16_io_data_out; // @[quant.scala 78:52]
  wire  unit_17_clock; // @[quant.scala 78:52]
  wire  unit_17_reset; // @[quant.scala 78:52]
  wire [7:0] unit_17_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_17_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_17_io_data_out; // @[quant.scala 78:52]
  wire  unit_18_clock; // @[quant.scala 78:52]
  wire  unit_18_reset; // @[quant.scala 78:52]
  wire [7:0] unit_18_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_18_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_18_io_data_out; // @[quant.scala 78:52]
  wire  unit_19_clock; // @[quant.scala 78:52]
  wire  unit_19_reset; // @[quant.scala 78:52]
  wire [7:0] unit_19_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_19_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_19_io_data_out; // @[quant.scala 78:52]
  wire  unit_20_clock; // @[quant.scala 78:52]
  wire  unit_20_reset; // @[quant.scala 78:52]
  wire [7:0] unit_20_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_20_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_20_io_data_out; // @[quant.scala 78:52]
  wire  unit_21_clock; // @[quant.scala 78:52]
  wire  unit_21_reset; // @[quant.scala 78:52]
  wire [7:0] unit_21_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_21_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_21_io_data_out; // @[quant.scala 78:52]
  wire  unit_22_clock; // @[quant.scala 78:52]
  wire  unit_22_reset; // @[quant.scala 78:52]
  wire [7:0] unit_22_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_22_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_22_io_data_out; // @[quant.scala 78:52]
  wire  unit_23_clock; // @[quant.scala 78:52]
  wire  unit_23_reset; // @[quant.scala 78:52]
  wire [7:0] unit_23_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_23_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_23_io_data_out; // @[quant.scala 78:52]
  wire  unit_24_clock; // @[quant.scala 78:52]
  wire  unit_24_reset; // @[quant.scala 78:52]
  wire [7:0] unit_24_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_24_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_24_io_data_out; // @[quant.scala 78:52]
  wire  unit_25_clock; // @[quant.scala 78:52]
  wire  unit_25_reset; // @[quant.scala 78:52]
  wire [7:0] unit_25_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_25_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_25_io_data_out; // @[quant.scala 78:52]
  wire  unit_26_clock; // @[quant.scala 78:52]
  wire  unit_26_reset; // @[quant.scala 78:52]
  wire [7:0] unit_26_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_26_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_26_io_data_out; // @[quant.scala 78:52]
  wire  unit_27_clock; // @[quant.scala 78:52]
  wire  unit_27_reset; // @[quant.scala 78:52]
  wire [7:0] unit_27_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_27_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_27_io_data_out; // @[quant.scala 78:52]
  wire  unit_28_clock; // @[quant.scala 78:52]
  wire  unit_28_reset; // @[quant.scala 78:52]
  wire [7:0] unit_28_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_28_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_28_io_data_out; // @[quant.scala 78:52]
  wire  unit_29_clock; // @[quant.scala 78:52]
  wire  unit_29_reset; // @[quant.scala 78:52]
  wire [7:0] unit_29_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_29_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_29_io_data_out; // @[quant.scala 78:52]
  wire  unit_30_clock; // @[quant.scala 78:52]
  wire  unit_30_reset; // @[quant.scala 78:52]
  wire [7:0] unit_30_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_30_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_30_io_data_out; // @[quant.scala 78:52]
  wire  unit_31_clock; // @[quant.scala 78:52]
  wire  unit_31_reset; // @[quant.scala 78:52]
  wire [7:0] unit_31_io_zero_point; // @[quant.scala 78:52]
  wire [7:0] unit_31_io_data_in; // @[quant.scala 78:52]
  wire [7:0] unit_31_io_data_out; // @[quant.scala 78:52]
  cal_sub_zero_point unit_0 ( // @[quant.scala 78:52]
    .clock(unit_0_clock),
    .reset(unit_0_reset),
    .io_zero_point(unit_0_io_zero_point),
    .io_data_in(unit_0_io_data_in),
    .io_data_out(unit_0_io_data_out)
  );
  cal_sub_zero_point unit_1 ( // @[quant.scala 78:52]
    .clock(unit_1_clock),
    .reset(unit_1_reset),
    .io_zero_point(unit_1_io_zero_point),
    .io_data_in(unit_1_io_data_in),
    .io_data_out(unit_1_io_data_out)
  );
  cal_sub_zero_point unit_2 ( // @[quant.scala 78:52]
    .clock(unit_2_clock),
    .reset(unit_2_reset),
    .io_zero_point(unit_2_io_zero_point),
    .io_data_in(unit_2_io_data_in),
    .io_data_out(unit_2_io_data_out)
  );
  cal_sub_zero_point unit_3 ( // @[quant.scala 78:52]
    .clock(unit_3_clock),
    .reset(unit_3_reset),
    .io_zero_point(unit_3_io_zero_point),
    .io_data_in(unit_3_io_data_in),
    .io_data_out(unit_3_io_data_out)
  );
  cal_sub_zero_point unit_4 ( // @[quant.scala 78:52]
    .clock(unit_4_clock),
    .reset(unit_4_reset),
    .io_zero_point(unit_4_io_zero_point),
    .io_data_in(unit_4_io_data_in),
    .io_data_out(unit_4_io_data_out)
  );
  cal_sub_zero_point unit_5 ( // @[quant.scala 78:52]
    .clock(unit_5_clock),
    .reset(unit_5_reset),
    .io_zero_point(unit_5_io_zero_point),
    .io_data_in(unit_5_io_data_in),
    .io_data_out(unit_5_io_data_out)
  );
  cal_sub_zero_point unit_6 ( // @[quant.scala 78:52]
    .clock(unit_6_clock),
    .reset(unit_6_reset),
    .io_zero_point(unit_6_io_zero_point),
    .io_data_in(unit_6_io_data_in),
    .io_data_out(unit_6_io_data_out)
  );
  cal_sub_zero_point unit_7 ( // @[quant.scala 78:52]
    .clock(unit_7_clock),
    .reset(unit_7_reset),
    .io_zero_point(unit_7_io_zero_point),
    .io_data_in(unit_7_io_data_in),
    .io_data_out(unit_7_io_data_out)
  );
  cal_sub_zero_point unit_8 ( // @[quant.scala 78:52]
    .clock(unit_8_clock),
    .reset(unit_8_reset),
    .io_zero_point(unit_8_io_zero_point),
    .io_data_in(unit_8_io_data_in),
    .io_data_out(unit_8_io_data_out)
  );
  cal_sub_zero_point unit_9 ( // @[quant.scala 78:52]
    .clock(unit_9_clock),
    .reset(unit_9_reset),
    .io_zero_point(unit_9_io_zero_point),
    .io_data_in(unit_9_io_data_in),
    .io_data_out(unit_9_io_data_out)
  );
  cal_sub_zero_point unit_10 ( // @[quant.scala 78:52]
    .clock(unit_10_clock),
    .reset(unit_10_reset),
    .io_zero_point(unit_10_io_zero_point),
    .io_data_in(unit_10_io_data_in),
    .io_data_out(unit_10_io_data_out)
  );
  cal_sub_zero_point unit_11 ( // @[quant.scala 78:52]
    .clock(unit_11_clock),
    .reset(unit_11_reset),
    .io_zero_point(unit_11_io_zero_point),
    .io_data_in(unit_11_io_data_in),
    .io_data_out(unit_11_io_data_out)
  );
  cal_sub_zero_point unit_12 ( // @[quant.scala 78:52]
    .clock(unit_12_clock),
    .reset(unit_12_reset),
    .io_zero_point(unit_12_io_zero_point),
    .io_data_in(unit_12_io_data_in),
    .io_data_out(unit_12_io_data_out)
  );
  cal_sub_zero_point unit_13 ( // @[quant.scala 78:52]
    .clock(unit_13_clock),
    .reset(unit_13_reset),
    .io_zero_point(unit_13_io_zero_point),
    .io_data_in(unit_13_io_data_in),
    .io_data_out(unit_13_io_data_out)
  );
  cal_sub_zero_point unit_14 ( // @[quant.scala 78:52]
    .clock(unit_14_clock),
    .reset(unit_14_reset),
    .io_zero_point(unit_14_io_zero_point),
    .io_data_in(unit_14_io_data_in),
    .io_data_out(unit_14_io_data_out)
  );
  cal_sub_zero_point unit_15 ( // @[quant.scala 78:52]
    .clock(unit_15_clock),
    .reset(unit_15_reset),
    .io_zero_point(unit_15_io_zero_point),
    .io_data_in(unit_15_io_data_in),
    .io_data_out(unit_15_io_data_out)
  );
  cal_sub_zero_point unit_16 ( // @[quant.scala 78:52]
    .clock(unit_16_clock),
    .reset(unit_16_reset),
    .io_zero_point(unit_16_io_zero_point),
    .io_data_in(unit_16_io_data_in),
    .io_data_out(unit_16_io_data_out)
  );
  cal_sub_zero_point unit_17 ( // @[quant.scala 78:52]
    .clock(unit_17_clock),
    .reset(unit_17_reset),
    .io_zero_point(unit_17_io_zero_point),
    .io_data_in(unit_17_io_data_in),
    .io_data_out(unit_17_io_data_out)
  );
  cal_sub_zero_point unit_18 ( // @[quant.scala 78:52]
    .clock(unit_18_clock),
    .reset(unit_18_reset),
    .io_zero_point(unit_18_io_zero_point),
    .io_data_in(unit_18_io_data_in),
    .io_data_out(unit_18_io_data_out)
  );
  cal_sub_zero_point unit_19 ( // @[quant.scala 78:52]
    .clock(unit_19_clock),
    .reset(unit_19_reset),
    .io_zero_point(unit_19_io_zero_point),
    .io_data_in(unit_19_io_data_in),
    .io_data_out(unit_19_io_data_out)
  );
  cal_sub_zero_point unit_20 ( // @[quant.scala 78:52]
    .clock(unit_20_clock),
    .reset(unit_20_reset),
    .io_zero_point(unit_20_io_zero_point),
    .io_data_in(unit_20_io_data_in),
    .io_data_out(unit_20_io_data_out)
  );
  cal_sub_zero_point unit_21 ( // @[quant.scala 78:52]
    .clock(unit_21_clock),
    .reset(unit_21_reset),
    .io_zero_point(unit_21_io_zero_point),
    .io_data_in(unit_21_io_data_in),
    .io_data_out(unit_21_io_data_out)
  );
  cal_sub_zero_point unit_22 ( // @[quant.scala 78:52]
    .clock(unit_22_clock),
    .reset(unit_22_reset),
    .io_zero_point(unit_22_io_zero_point),
    .io_data_in(unit_22_io_data_in),
    .io_data_out(unit_22_io_data_out)
  );
  cal_sub_zero_point unit_23 ( // @[quant.scala 78:52]
    .clock(unit_23_clock),
    .reset(unit_23_reset),
    .io_zero_point(unit_23_io_zero_point),
    .io_data_in(unit_23_io_data_in),
    .io_data_out(unit_23_io_data_out)
  );
  cal_sub_zero_point unit_24 ( // @[quant.scala 78:52]
    .clock(unit_24_clock),
    .reset(unit_24_reset),
    .io_zero_point(unit_24_io_zero_point),
    .io_data_in(unit_24_io_data_in),
    .io_data_out(unit_24_io_data_out)
  );
  cal_sub_zero_point unit_25 ( // @[quant.scala 78:52]
    .clock(unit_25_clock),
    .reset(unit_25_reset),
    .io_zero_point(unit_25_io_zero_point),
    .io_data_in(unit_25_io_data_in),
    .io_data_out(unit_25_io_data_out)
  );
  cal_sub_zero_point unit_26 ( // @[quant.scala 78:52]
    .clock(unit_26_clock),
    .reset(unit_26_reset),
    .io_zero_point(unit_26_io_zero_point),
    .io_data_in(unit_26_io_data_in),
    .io_data_out(unit_26_io_data_out)
  );
  cal_sub_zero_point unit_27 ( // @[quant.scala 78:52]
    .clock(unit_27_clock),
    .reset(unit_27_reset),
    .io_zero_point(unit_27_io_zero_point),
    .io_data_in(unit_27_io_data_in),
    .io_data_out(unit_27_io_data_out)
  );
  cal_sub_zero_point unit_28 ( // @[quant.scala 78:52]
    .clock(unit_28_clock),
    .reset(unit_28_reset),
    .io_zero_point(unit_28_io_zero_point),
    .io_data_in(unit_28_io_data_in),
    .io_data_out(unit_28_io_data_out)
  );
  cal_sub_zero_point unit_29 ( // @[quant.scala 78:52]
    .clock(unit_29_clock),
    .reset(unit_29_reset),
    .io_zero_point(unit_29_io_zero_point),
    .io_data_in(unit_29_io_data_in),
    .io_data_out(unit_29_io_data_out)
  );
  cal_sub_zero_point unit_30 ( // @[quant.scala 78:52]
    .clock(unit_30_clock),
    .reset(unit_30_reset),
    .io_zero_point(unit_30_io_zero_point),
    .io_data_in(unit_30_io_data_in),
    .io_data_out(unit_30_io_data_out)
  );
  cal_sub_zero_point unit_31 ( // @[quant.scala 78:52]
    .clock(unit_31_clock),
    .reset(unit_31_reset),
    .io_zero_point(unit_31_io_zero_point),
    .io_data_in(unit_31_io_data_in),
    .io_data_out(unit_31_io_data_out)
  );
  assign io_data_out_0 = unit_0_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_1 = unit_1_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_2 = unit_2_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_3 = unit_3_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_4 = unit_4_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_5 = unit_5_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_6 = unit_6_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_7 = unit_7_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_8 = unit_8_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_9 = unit_9_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_10 = unit_10_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_11 = unit_11_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_12 = unit_12_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_13 = unit_13_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_14 = unit_14_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_15 = unit_15_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_16 = unit_16_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_17 = unit_17_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_18 = unit_18_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_19 = unit_19_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_20 = unit_20_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_21 = unit_21_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_22 = unit_22_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_23 = unit_23_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_24 = unit_24_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_25 = unit_25_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_26 = unit_26_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_27 = unit_27_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_28 = unit_28_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_29 = unit_29_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_30 = unit_30_io_data_out; // @[quant.scala 82:24]
  assign io_data_out_31 = unit_31_io_data_out; // @[quant.scala 82:24]
  assign unit_0_clock = clock;
  assign unit_0_reset = reset;
  assign unit_0_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_0_io_data_in = io_data_in_0; // @[quant.scala 81:28]
  assign unit_1_clock = clock;
  assign unit_1_reset = reset;
  assign unit_1_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_1_io_data_in = io_data_in_1; // @[quant.scala 81:28]
  assign unit_2_clock = clock;
  assign unit_2_reset = reset;
  assign unit_2_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_2_io_data_in = io_data_in_2; // @[quant.scala 81:28]
  assign unit_3_clock = clock;
  assign unit_3_reset = reset;
  assign unit_3_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_3_io_data_in = io_data_in_3; // @[quant.scala 81:28]
  assign unit_4_clock = clock;
  assign unit_4_reset = reset;
  assign unit_4_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_4_io_data_in = io_data_in_4; // @[quant.scala 81:28]
  assign unit_5_clock = clock;
  assign unit_5_reset = reset;
  assign unit_5_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_5_io_data_in = io_data_in_5; // @[quant.scala 81:28]
  assign unit_6_clock = clock;
  assign unit_6_reset = reset;
  assign unit_6_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_6_io_data_in = io_data_in_6; // @[quant.scala 81:28]
  assign unit_7_clock = clock;
  assign unit_7_reset = reset;
  assign unit_7_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_7_io_data_in = io_data_in_7; // @[quant.scala 81:28]
  assign unit_8_clock = clock;
  assign unit_8_reset = reset;
  assign unit_8_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_8_io_data_in = io_data_in_8; // @[quant.scala 81:28]
  assign unit_9_clock = clock;
  assign unit_9_reset = reset;
  assign unit_9_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_9_io_data_in = io_data_in_9; // @[quant.scala 81:28]
  assign unit_10_clock = clock;
  assign unit_10_reset = reset;
  assign unit_10_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_10_io_data_in = io_data_in_10; // @[quant.scala 81:28]
  assign unit_11_clock = clock;
  assign unit_11_reset = reset;
  assign unit_11_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_11_io_data_in = io_data_in_11; // @[quant.scala 81:28]
  assign unit_12_clock = clock;
  assign unit_12_reset = reset;
  assign unit_12_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_12_io_data_in = io_data_in_12; // @[quant.scala 81:28]
  assign unit_13_clock = clock;
  assign unit_13_reset = reset;
  assign unit_13_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_13_io_data_in = io_data_in_13; // @[quant.scala 81:28]
  assign unit_14_clock = clock;
  assign unit_14_reset = reset;
  assign unit_14_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_14_io_data_in = io_data_in_14; // @[quant.scala 81:28]
  assign unit_15_clock = clock;
  assign unit_15_reset = reset;
  assign unit_15_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_15_io_data_in = io_data_in_15; // @[quant.scala 81:28]
  assign unit_16_clock = clock;
  assign unit_16_reset = reset;
  assign unit_16_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_16_io_data_in = io_data_in_16; // @[quant.scala 81:28]
  assign unit_17_clock = clock;
  assign unit_17_reset = reset;
  assign unit_17_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_17_io_data_in = io_data_in_17; // @[quant.scala 81:28]
  assign unit_18_clock = clock;
  assign unit_18_reset = reset;
  assign unit_18_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_18_io_data_in = io_data_in_18; // @[quant.scala 81:28]
  assign unit_19_clock = clock;
  assign unit_19_reset = reset;
  assign unit_19_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_19_io_data_in = io_data_in_19; // @[quant.scala 81:28]
  assign unit_20_clock = clock;
  assign unit_20_reset = reset;
  assign unit_20_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_20_io_data_in = io_data_in_20; // @[quant.scala 81:28]
  assign unit_21_clock = clock;
  assign unit_21_reset = reset;
  assign unit_21_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_21_io_data_in = io_data_in_21; // @[quant.scala 81:28]
  assign unit_22_clock = clock;
  assign unit_22_reset = reset;
  assign unit_22_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_22_io_data_in = io_data_in_22; // @[quant.scala 81:28]
  assign unit_23_clock = clock;
  assign unit_23_reset = reset;
  assign unit_23_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_23_io_data_in = io_data_in_23; // @[quant.scala 81:28]
  assign unit_24_clock = clock;
  assign unit_24_reset = reset;
  assign unit_24_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_24_io_data_in = io_data_in_24; // @[quant.scala 81:28]
  assign unit_25_clock = clock;
  assign unit_25_reset = reset;
  assign unit_25_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_25_io_data_in = io_data_in_25; // @[quant.scala 81:28]
  assign unit_26_clock = clock;
  assign unit_26_reset = reset;
  assign unit_26_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_26_io_data_in = io_data_in_26; // @[quant.scala 81:28]
  assign unit_27_clock = clock;
  assign unit_27_reset = reset;
  assign unit_27_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_27_io_data_in = io_data_in_27; // @[quant.scala 81:28]
  assign unit_28_clock = clock;
  assign unit_28_reset = reset;
  assign unit_28_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_28_io_data_in = io_data_in_28; // @[quant.scala 81:28]
  assign unit_29_clock = clock;
  assign unit_29_reset = reset;
  assign unit_29_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_29_io_data_in = io_data_in_29; // @[quant.scala 81:28]
  assign unit_30_clock = clock;
  assign unit_30_reset = reset;
  assign unit_30_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_30_io_data_in = io_data_in_30; // @[quant.scala 81:28]
  assign unit_31_clock = clock;
  assign unit_31_reset = reset;
  assign unit_31_io_zero_point = io_zero_point; // @[quant.scala 80:31]
  assign unit_31_io_data_in = io_data_in_31; // @[quant.scala 81:28]
endmodule
module linebuf_unit_extend(
  input         clock,
  input         reset,
  input  [15:0] io_i,
  output [15:0] io_o,
  input         io_s_mod,
  input         io_line_extend_en,
  input  [2:0]  io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] reg_temp0; // @[LineBuffer.scala 99:28]
  reg [7:0] reg_temp1; // @[LineBuffer.scala 100:28]
  reg [7:0] reg_temp2; // @[LineBuffer.scala 101:28]
  reg [7:0] line_shift_1_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_39; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_40; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_41; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_42; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_43; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_44; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_45; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_46; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_47; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_48; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_49; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_50; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_51; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_52; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_53; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_54; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_55; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_56; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_57; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_58; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_59; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_60; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_61; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_62; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_63; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_64; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_65; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_66; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_67; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_68; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_69; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_70; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_71; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_72; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_73; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_74; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_75; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_76; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_77; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_78; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_39; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_40; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_41; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_42; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_43; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_44; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_45; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_46; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_47; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_48; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_49; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_50; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_51; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_52; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_53; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_54; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_55; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_56; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_57; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_58; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_59; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_60; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_61; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_62; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_63; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_64; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_65; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_66; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_67; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_68; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_69; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_70; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_71; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_72; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_73; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_74; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_75; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_76; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_77; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_78; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_79; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_80; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_81; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_82; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_83; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_84; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_85; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_86; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_87; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_88; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_89; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_90; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_91; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_92; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_93; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_94; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_95; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_96; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_97; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_98; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_99; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_100; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_101; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_102; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_103; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_104; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_105; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_106; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_107; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_108; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_109; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_110; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_111; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_112; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_113; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_114; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_115; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_116; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_117; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_118; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_119; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_120; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_121; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_122; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_123; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_124; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_125; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_126; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_127; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_128; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_129; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_130; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_131; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_132; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_133; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_134; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_135; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_136; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_137; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_138; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_139; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_140; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_141; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_142; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_143; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_144; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_145; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_146; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_147; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_148; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_149; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_150; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_151; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_152; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_153; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_154; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_155; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_156; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_157; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5_r_158; // @[Reg.scala 35:20]
  reg [7:0] line_shift_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_39; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_40; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_41; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_42; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_43; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_44; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_45; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_46; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_47; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_48; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_49; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_50; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_51; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_52; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_53; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_54; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_55; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_56; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_57; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_58; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_59; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_60; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_61; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_62; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_63; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_64; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_65; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_66; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_67; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_68; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_69; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_70; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_71; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_72; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_73; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_74; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_75; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_76; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_77; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14_r_78; // @[Reg.scala 35:20]
  reg [7:0] line_shift_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_19; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_20; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_21; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_22; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_23; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_24; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_25; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_26; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_27; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_28; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_29; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_30; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_31; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_32; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_33; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_34; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_35; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_36; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_37; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_38; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_39; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_40; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_41; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_42; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_43; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_44; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_45; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_46; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_47; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_48; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_49; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_50; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_51; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_52; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_53; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_54; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_55; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_56; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_57; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_58; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_59; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_60; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_61; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_62; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_63; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_64; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_65; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_66; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_67; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_68; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_69; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_70; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_71; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_72; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_73; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_74; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_75; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_76; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_77; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_78; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_79; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_80; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_81; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_82; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_83; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_84; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_85; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_86; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_87; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_88; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_89; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_90; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_91; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_92; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_93; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_94; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_95; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_96; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_97; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_98; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_99; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_100; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_101; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_102; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_103; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_104; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_105; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_106; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_107; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_108; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_109; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_110; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_111; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_112; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_113; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_114; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_115; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_116; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_117; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_118; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_119; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_120; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_121; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_122; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_123; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_124; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_125; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_126; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_127; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_128; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_129; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_130; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_131; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_132; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_133; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_134; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_135; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_136; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_137; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_138; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_139; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_140; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_141; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_142; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_143; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_144; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_145; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_146; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_147; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_148; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_149; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_150; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_151; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_152; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_153; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_154; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_155; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_156; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_157; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15_r_158; // @[Reg.scala 35:20]
  reg [7:0] line_shift_15; // @[Reg.scala 35:20]
  wire [7:0] _temp_out_0_T_1 = 3'h0 == io_sel ? line_shift_1 : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_0_T_3 = 3'h1 == io_sel ? line_shift_2 : _temp_out_0_T_1; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_0_T_5 = 3'h2 == io_sel ? line_shift_3 : _temp_out_0_T_3; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_0_T_7 = 3'h3 == io_sel ? line_shift_4 : _temp_out_0_T_5; // @[Mux.scala 81:58]
  wire [7:0] temp_out_0 = 3'h4 == io_sel ? line_shift_5 : _temp_out_0_T_7; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_1_T_1 = 3'h0 == io_sel ? line_shift_11 : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_1_T_3 = 3'h1 == io_sel ? line_shift_12 : _temp_out_1_T_1; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_1_T_5 = 3'h2 == io_sel ? line_shift_13 : _temp_out_1_T_3; // @[Mux.scala 81:58]
  wire [7:0] _temp_out_1_T_7 = 3'h3 == io_sel ? line_shift_14 : _temp_out_1_T_5; // @[Mux.scala 81:58]
  wire [7:0] temp_out_1 = 3'h4 == io_sel ? line_shift_15 : _temp_out_1_T_7; // @[Mux.scala 81:58]
  assign io_o = {temp_out_1,temp_out_0}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[LineBuffer.scala 99:28]
      reg_temp0 <= 8'h0; // @[LineBuffer.scala 99:28]
    end else begin
      reg_temp0 <= io_i[7:0]; // @[LineBuffer.scala 102:15]
    end
    if (reset) begin // @[LineBuffer.scala 100:28]
      reg_temp1 <= 8'h0; // @[LineBuffer.scala 100:28]
    end else begin
      reg_temp1 <= io_i[15:8]; // @[LineBuffer.scala 103:15]
    end
    if (reset) begin // @[LineBuffer.scala 101:28]
      reg_temp2 <= 8'h0; // @[LineBuffer.scala 101:28]
    end else begin
      reg_temp2 <= reg_temp0; // @[LineBuffer.scala 104:15]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_s_mod) begin // @[LineBuffer.scala 106:36]
      line_shift_1_r <= reg_temp0;
    end else begin
      line_shift_1_r <= reg_temp2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_1 <= line_shift_1_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_2 <= line_shift_1_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_3 <= line_shift_1_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_4 <= line_shift_1_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_5 <= line_shift_1_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_6 <= line_shift_1_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_7 <= line_shift_1_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_8 <= line_shift_1_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_9 <= line_shift_1_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_10 <= line_shift_1_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_11 <= line_shift_1_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_12 <= line_shift_1_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_13 <= line_shift_1_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_14 <= line_shift_1_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_15 <= line_shift_1_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_16 <= line_shift_1_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_17 <= line_shift_1_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1_r_18 <= line_shift_1_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_1 <= line_shift_1_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r <= line_shift_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_1 <= line_shift_2_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_2 <= line_shift_2_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_3 <= line_shift_2_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_4 <= line_shift_2_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_5 <= line_shift_2_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_6 <= line_shift_2_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_7 <= line_shift_2_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_8 <= line_shift_2_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_9 <= line_shift_2_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_10 <= line_shift_2_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_11 <= line_shift_2_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_12 <= line_shift_2_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_13 <= line_shift_2_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_14 <= line_shift_2_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_15 <= line_shift_2_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_16 <= line_shift_2_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_17 <= line_shift_2_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2_r_18 <= line_shift_2_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_2 <= line_shift_2_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r <= line_shift_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_1 <= line_shift_3_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_2 <= line_shift_3_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_3 <= line_shift_3_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_4 <= line_shift_3_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_5 <= line_shift_3_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_6 <= line_shift_3_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_7 <= line_shift_3_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_8 <= line_shift_3_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_9 <= line_shift_3_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_10 <= line_shift_3_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_11 <= line_shift_3_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_12 <= line_shift_3_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_13 <= line_shift_3_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_14 <= line_shift_3_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_15 <= line_shift_3_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_16 <= line_shift_3_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_17 <= line_shift_3_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_18 <= line_shift_3_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_19 <= line_shift_3_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_20 <= line_shift_3_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_21 <= line_shift_3_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_22 <= line_shift_3_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_23 <= line_shift_3_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_24 <= line_shift_3_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_25 <= line_shift_3_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_26 <= line_shift_3_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_27 <= line_shift_3_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_28 <= line_shift_3_r_27;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_29 <= line_shift_3_r_28;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_30 <= line_shift_3_r_29;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_31 <= line_shift_3_r_30;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_32 <= line_shift_3_r_31;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_33 <= line_shift_3_r_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_34 <= line_shift_3_r_33;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_35 <= line_shift_3_r_34;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_36 <= line_shift_3_r_35;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_37 <= line_shift_3_r_36;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3_r_38 <= line_shift_3_r_37;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_3 <= line_shift_3_r_38;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r <= line_shift_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_1 <= line_shift_4_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_2 <= line_shift_4_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_3 <= line_shift_4_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_4 <= line_shift_4_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_5 <= line_shift_4_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_6 <= line_shift_4_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_7 <= line_shift_4_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_8 <= line_shift_4_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_9 <= line_shift_4_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_10 <= line_shift_4_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_11 <= line_shift_4_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_12 <= line_shift_4_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_13 <= line_shift_4_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_14 <= line_shift_4_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_15 <= line_shift_4_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_16 <= line_shift_4_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_17 <= line_shift_4_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_18 <= line_shift_4_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_19 <= line_shift_4_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_20 <= line_shift_4_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_21 <= line_shift_4_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_22 <= line_shift_4_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_23 <= line_shift_4_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_24 <= line_shift_4_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_25 <= line_shift_4_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_26 <= line_shift_4_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_27 <= line_shift_4_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_28 <= line_shift_4_r_27;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_29 <= line_shift_4_r_28;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_30 <= line_shift_4_r_29;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_31 <= line_shift_4_r_30;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_32 <= line_shift_4_r_31;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_33 <= line_shift_4_r_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_34 <= line_shift_4_r_33;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_35 <= line_shift_4_r_34;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_36 <= line_shift_4_r_35;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_37 <= line_shift_4_r_36;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_38 <= line_shift_4_r_37;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_39 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_39 <= line_shift_4_r_38;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_40 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_40 <= line_shift_4_r_39;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_41 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_41 <= line_shift_4_r_40;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_42 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_42 <= line_shift_4_r_41;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_43 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_43 <= line_shift_4_r_42;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_44 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_44 <= line_shift_4_r_43;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_45 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_45 <= line_shift_4_r_44;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_46 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_46 <= line_shift_4_r_45;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_47 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_47 <= line_shift_4_r_46;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_48 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_48 <= line_shift_4_r_47;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_49 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_49 <= line_shift_4_r_48;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_50 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_50 <= line_shift_4_r_49;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_51 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_51 <= line_shift_4_r_50;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_52 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_52 <= line_shift_4_r_51;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_53 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_53 <= line_shift_4_r_52;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_54 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_54 <= line_shift_4_r_53;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_55 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_55 <= line_shift_4_r_54;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_56 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_56 <= line_shift_4_r_55;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_57 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_57 <= line_shift_4_r_56;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_58 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_58 <= line_shift_4_r_57;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_59 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_59 <= line_shift_4_r_58;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_60 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_60 <= line_shift_4_r_59;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_61 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_61 <= line_shift_4_r_60;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_62 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_62 <= line_shift_4_r_61;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_63 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_63 <= line_shift_4_r_62;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_64 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_64 <= line_shift_4_r_63;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_65 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_65 <= line_shift_4_r_64;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_66 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_66 <= line_shift_4_r_65;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_67 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_67 <= line_shift_4_r_66;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_68 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_68 <= line_shift_4_r_67;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_69 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_69 <= line_shift_4_r_68;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_70 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_70 <= line_shift_4_r_69;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_71 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_71 <= line_shift_4_r_70;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_72 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_72 <= line_shift_4_r_71;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_73 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_73 <= line_shift_4_r_72;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_74 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_74 <= line_shift_4_r_73;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_75 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_75 <= line_shift_4_r_74;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_76 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_76 <= line_shift_4_r_75;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_77 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_77 <= line_shift_4_r_76;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_78 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4_r_78 <= line_shift_4_r_77;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_4 <= line_shift_4_r_78;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r <= line_shift_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_1 <= line_shift_5_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_2 <= line_shift_5_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_3 <= line_shift_5_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_4 <= line_shift_5_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_5 <= line_shift_5_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_6 <= line_shift_5_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_7 <= line_shift_5_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_8 <= line_shift_5_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_9 <= line_shift_5_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_10 <= line_shift_5_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_11 <= line_shift_5_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_12 <= line_shift_5_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_13 <= line_shift_5_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_14 <= line_shift_5_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_15 <= line_shift_5_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_16 <= line_shift_5_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_17 <= line_shift_5_r_16;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_18 <= line_shift_5_r_17;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_19 <= line_shift_5_r_18;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_20 <= line_shift_5_r_19;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_21 <= line_shift_5_r_20;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_22 <= line_shift_5_r_21;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_23 <= line_shift_5_r_22;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_24 <= line_shift_5_r_23;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_25 <= line_shift_5_r_24;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_26 <= line_shift_5_r_25;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_27 <= line_shift_5_r_26;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_28 <= line_shift_5_r_27;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_29 <= line_shift_5_r_28;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_30 <= line_shift_5_r_29;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_31 <= line_shift_5_r_30;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_32 <= line_shift_5_r_31;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_33 <= line_shift_5_r_32;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_34 <= line_shift_5_r_33;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_35 <= line_shift_5_r_34;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_36 <= line_shift_5_r_35;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_37 <= line_shift_5_r_36;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_38 <= line_shift_5_r_37;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_39 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_39 <= line_shift_5_r_38;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_40 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_40 <= line_shift_5_r_39;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_41 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_41 <= line_shift_5_r_40;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_42 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_42 <= line_shift_5_r_41;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_43 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_43 <= line_shift_5_r_42;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_44 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_44 <= line_shift_5_r_43;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_45 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_45 <= line_shift_5_r_44;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_46 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_46 <= line_shift_5_r_45;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_47 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_47 <= line_shift_5_r_46;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_48 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_48 <= line_shift_5_r_47;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_49 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_49 <= line_shift_5_r_48;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_50 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_50 <= line_shift_5_r_49;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_51 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_51 <= line_shift_5_r_50;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_52 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_52 <= line_shift_5_r_51;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_53 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_53 <= line_shift_5_r_52;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_54 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_54 <= line_shift_5_r_53;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_55 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_55 <= line_shift_5_r_54;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_56 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_56 <= line_shift_5_r_55;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_57 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_57 <= line_shift_5_r_56;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_58 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_58 <= line_shift_5_r_57;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_59 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_59 <= line_shift_5_r_58;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_60 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_60 <= line_shift_5_r_59;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_61 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_61 <= line_shift_5_r_60;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_62 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_62 <= line_shift_5_r_61;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_63 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_63 <= line_shift_5_r_62;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_64 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_64 <= line_shift_5_r_63;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_65 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_65 <= line_shift_5_r_64;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_66 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_66 <= line_shift_5_r_65;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_67 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_67 <= line_shift_5_r_66;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_68 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_68 <= line_shift_5_r_67;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_69 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_69 <= line_shift_5_r_68;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_70 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_70 <= line_shift_5_r_69;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_71 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_71 <= line_shift_5_r_70;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_72 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_72 <= line_shift_5_r_71;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_73 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_73 <= line_shift_5_r_72;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_74 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_74 <= line_shift_5_r_73;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_75 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_75 <= line_shift_5_r_74;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_76 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_76 <= line_shift_5_r_75;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_77 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_77 <= line_shift_5_r_76;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_78 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_78 <= line_shift_5_r_77;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_79 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_79 <= line_shift_5_r_78;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_80 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_80 <= line_shift_5_r_79;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_81 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_81 <= line_shift_5_r_80;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_82 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_82 <= line_shift_5_r_81;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_83 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_83 <= line_shift_5_r_82;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_84 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_84 <= line_shift_5_r_83;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_85 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_85 <= line_shift_5_r_84;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_86 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_86 <= line_shift_5_r_85;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_87 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_87 <= line_shift_5_r_86;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_88 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_88 <= line_shift_5_r_87;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_89 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_89 <= line_shift_5_r_88;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_90 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_90 <= line_shift_5_r_89;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_91 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_91 <= line_shift_5_r_90;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_92 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_92 <= line_shift_5_r_91;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_93 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_93 <= line_shift_5_r_92;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_94 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_94 <= line_shift_5_r_93;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_95 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_95 <= line_shift_5_r_94;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_96 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_96 <= line_shift_5_r_95;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_97 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_97 <= line_shift_5_r_96;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_98 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_98 <= line_shift_5_r_97;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_99 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_99 <= line_shift_5_r_98;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_100 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_100 <= line_shift_5_r_99;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_101 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_101 <= line_shift_5_r_100;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_102 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_102 <= line_shift_5_r_101;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_103 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_103 <= line_shift_5_r_102;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_104 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_104 <= line_shift_5_r_103;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_105 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_105 <= line_shift_5_r_104;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_106 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_106 <= line_shift_5_r_105;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_107 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_107 <= line_shift_5_r_106;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_108 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_108 <= line_shift_5_r_107;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_109 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_109 <= line_shift_5_r_108;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_110 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_110 <= line_shift_5_r_109;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_111 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_111 <= line_shift_5_r_110;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_112 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_112 <= line_shift_5_r_111;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_113 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_113 <= line_shift_5_r_112;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_114 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_114 <= line_shift_5_r_113;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_115 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_115 <= line_shift_5_r_114;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_116 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_116 <= line_shift_5_r_115;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_117 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_117 <= line_shift_5_r_116;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_118 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_118 <= line_shift_5_r_117;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_119 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_119 <= line_shift_5_r_118;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_120 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_120 <= line_shift_5_r_119;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_121 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_121 <= line_shift_5_r_120;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_122 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_122 <= line_shift_5_r_121;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_123 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_123 <= line_shift_5_r_122;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_124 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_124 <= line_shift_5_r_123;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_125 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_125 <= line_shift_5_r_124;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_126 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_126 <= line_shift_5_r_125;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_127 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_127 <= line_shift_5_r_126;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_128 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_128 <= line_shift_5_r_127;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_129 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_129 <= line_shift_5_r_128;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_130 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_130 <= line_shift_5_r_129;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_131 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_131 <= line_shift_5_r_130;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_132 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_132 <= line_shift_5_r_131;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_133 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_133 <= line_shift_5_r_132;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_134 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_134 <= line_shift_5_r_133;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_135 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_135 <= line_shift_5_r_134;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_136 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_136 <= line_shift_5_r_135;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_137 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_137 <= line_shift_5_r_136;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_138 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_138 <= line_shift_5_r_137;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_139 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_139 <= line_shift_5_r_138;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_140 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_140 <= line_shift_5_r_139;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_141 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_141 <= line_shift_5_r_140;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_142 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_142 <= line_shift_5_r_141;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_143 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_143 <= line_shift_5_r_142;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_144 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_144 <= line_shift_5_r_143;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_145 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_145 <= line_shift_5_r_144;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_146 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_146 <= line_shift_5_r_145;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_147 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_147 <= line_shift_5_r_146;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_148 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_148 <= line_shift_5_r_147;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_149 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_149 <= line_shift_5_r_148;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_150 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_150 <= line_shift_5_r_149;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_151 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_151 <= line_shift_5_r_150;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_152 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_152 <= line_shift_5_r_151;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_153 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_153 <= line_shift_5_r_152;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_154 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_154 <= line_shift_5_r_153;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_155 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_155 <= line_shift_5_r_154;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_156 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_156 <= line_shift_5_r_155;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_157 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_157 <= line_shift_5_r_156;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5_r_158 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5_r_158 <= line_shift_5_r_157;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_5 <= 8'h0; // @[Reg.scala 35:20]
    end else begin
      line_shift_5 <= line_shift_5_r_158;
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r <= reg_temp1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_1 <= line_shift_11_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_2 <= line_shift_11_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_3 <= line_shift_11_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_4 <= line_shift_11_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_5 <= line_shift_11_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_6 <= line_shift_11_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_7 <= line_shift_11_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_8 <= line_shift_11_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_9 <= line_shift_11_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_10 <= line_shift_11_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_11 <= line_shift_11_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_12 <= line_shift_11_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_13 <= line_shift_11_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_14 <= line_shift_11_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_15 <= line_shift_11_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_16 <= line_shift_11_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_17 <= line_shift_11_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11_r_18 <= line_shift_11_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_11 <= line_shift_11_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r <= line_shift_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_1 <= line_shift_12_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_2 <= line_shift_12_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_3 <= line_shift_12_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_4 <= line_shift_12_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_5 <= line_shift_12_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_6 <= line_shift_12_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_7 <= line_shift_12_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_8 <= line_shift_12_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_9 <= line_shift_12_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_10 <= line_shift_12_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_11 <= line_shift_12_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_12 <= line_shift_12_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_13 <= line_shift_12_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_14 <= line_shift_12_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_15 <= line_shift_12_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_16 <= line_shift_12_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_17 <= line_shift_12_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12_r_18 <= line_shift_12_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_12 <= line_shift_12_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r <= line_shift_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_1 <= line_shift_13_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_2 <= line_shift_13_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_3 <= line_shift_13_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_4 <= line_shift_13_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_5 <= line_shift_13_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_6 <= line_shift_13_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_7 <= line_shift_13_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_8 <= line_shift_13_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_9 <= line_shift_13_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_10 <= line_shift_13_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_11 <= line_shift_13_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_12 <= line_shift_13_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_13 <= line_shift_13_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_14 <= line_shift_13_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_15 <= line_shift_13_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_16 <= line_shift_13_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_17 <= line_shift_13_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_18 <= line_shift_13_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_19 <= line_shift_13_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_20 <= line_shift_13_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_21 <= line_shift_13_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_22 <= line_shift_13_r_21; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_23 <= line_shift_13_r_22; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_24 <= line_shift_13_r_23; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_25 <= line_shift_13_r_24; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_26 <= line_shift_13_r_25; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_27 <= line_shift_13_r_26; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_28 <= line_shift_13_r_27; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_29 <= line_shift_13_r_28; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_30 <= line_shift_13_r_29; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_31 <= line_shift_13_r_30; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_32 <= line_shift_13_r_31; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_33 <= line_shift_13_r_32; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_34 <= line_shift_13_r_33; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_35 <= line_shift_13_r_34; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_36 <= line_shift_13_r_35; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_37 <= line_shift_13_r_36; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13_r_38 <= line_shift_13_r_37; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_13 <= line_shift_13_r_38; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r <= line_shift_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_1 <= line_shift_14_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_2 <= line_shift_14_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_3 <= line_shift_14_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_4 <= line_shift_14_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_5 <= line_shift_14_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_6 <= line_shift_14_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_7 <= line_shift_14_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_8 <= line_shift_14_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_9 <= line_shift_14_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_10 <= line_shift_14_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_11 <= line_shift_14_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_12 <= line_shift_14_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_13 <= line_shift_14_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_14 <= line_shift_14_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_15 <= line_shift_14_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_16 <= line_shift_14_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_17 <= line_shift_14_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_18 <= line_shift_14_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_19 <= line_shift_14_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_20 <= line_shift_14_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_21 <= line_shift_14_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_22 <= line_shift_14_r_21; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_23 <= line_shift_14_r_22; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_24 <= line_shift_14_r_23; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_25 <= line_shift_14_r_24; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_26 <= line_shift_14_r_25; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_27 <= line_shift_14_r_26; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_28 <= line_shift_14_r_27; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_29 <= line_shift_14_r_28; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_30 <= line_shift_14_r_29; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_31 <= line_shift_14_r_30; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_32 <= line_shift_14_r_31; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_33 <= line_shift_14_r_32; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_34 <= line_shift_14_r_33; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_35 <= line_shift_14_r_34; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_36 <= line_shift_14_r_35; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_37 <= line_shift_14_r_36; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_38 <= line_shift_14_r_37; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_39 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_39 <= line_shift_14_r_38; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_40 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_40 <= line_shift_14_r_39; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_41 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_41 <= line_shift_14_r_40; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_42 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_42 <= line_shift_14_r_41; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_43 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_43 <= line_shift_14_r_42; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_44 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_44 <= line_shift_14_r_43; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_45 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_45 <= line_shift_14_r_44; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_46 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_46 <= line_shift_14_r_45; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_47 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_47 <= line_shift_14_r_46; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_48 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_48 <= line_shift_14_r_47; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_49 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_49 <= line_shift_14_r_48; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_50 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_50 <= line_shift_14_r_49; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_51 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_51 <= line_shift_14_r_50; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_52 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_52 <= line_shift_14_r_51; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_53 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_53 <= line_shift_14_r_52; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_54 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_54 <= line_shift_14_r_53; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_55 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_55 <= line_shift_14_r_54; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_56 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_56 <= line_shift_14_r_55; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_57 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_57 <= line_shift_14_r_56; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_58 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_58 <= line_shift_14_r_57; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_59 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_59 <= line_shift_14_r_58; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_60 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_60 <= line_shift_14_r_59; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_61 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_61 <= line_shift_14_r_60; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_62 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_62 <= line_shift_14_r_61; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_63 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_63 <= line_shift_14_r_62; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_64 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_64 <= line_shift_14_r_63; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_65 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_65 <= line_shift_14_r_64; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_66 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_66 <= line_shift_14_r_65; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_67 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_67 <= line_shift_14_r_66; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_68 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_68 <= line_shift_14_r_67; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_69 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_69 <= line_shift_14_r_68; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_70 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_70 <= line_shift_14_r_69; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_71 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_71 <= line_shift_14_r_70; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_72 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_72 <= line_shift_14_r_71; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_73 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_73 <= line_shift_14_r_72; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_74 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_74 <= line_shift_14_r_73; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_75 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_75 <= line_shift_14_r_74; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_76 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_76 <= line_shift_14_r_75; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_77 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_77 <= line_shift_14_r_76; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14_r_78 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14_r_78 <= line_shift_14_r_77; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_14 <= line_shift_14_r_78; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r <= line_shift_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_1 <= line_shift_15_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_2 <= line_shift_15_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_3 <= line_shift_15_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_4 <= line_shift_15_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_5 <= line_shift_15_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_6 <= line_shift_15_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_7 <= line_shift_15_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_8 <= line_shift_15_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_9 <= line_shift_15_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_10 <= line_shift_15_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_11 <= line_shift_15_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_12 <= line_shift_15_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_13 <= line_shift_15_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_14 <= line_shift_15_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_15 <= line_shift_15_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_16 <= line_shift_15_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_17 <= line_shift_15_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_18 <= line_shift_15_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_19 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_19 <= line_shift_15_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_20 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_20 <= line_shift_15_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_21 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_21 <= line_shift_15_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_22 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_22 <= line_shift_15_r_21; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_23 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_23 <= line_shift_15_r_22; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_24 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_24 <= line_shift_15_r_23; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_25 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_25 <= line_shift_15_r_24; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_26 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_26 <= line_shift_15_r_25; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_27 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_27 <= line_shift_15_r_26; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_28 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_28 <= line_shift_15_r_27; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_29 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_29 <= line_shift_15_r_28; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_30 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_30 <= line_shift_15_r_29; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_31 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_31 <= line_shift_15_r_30; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_32 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_32 <= line_shift_15_r_31; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_33 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_33 <= line_shift_15_r_32; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_34 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_34 <= line_shift_15_r_33; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_35 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_35 <= line_shift_15_r_34; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_36 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_36 <= line_shift_15_r_35; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_37 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_37 <= line_shift_15_r_36; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_38 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_38 <= line_shift_15_r_37; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_39 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_39 <= line_shift_15_r_38; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_40 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_40 <= line_shift_15_r_39; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_41 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_41 <= line_shift_15_r_40; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_42 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_42 <= line_shift_15_r_41; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_43 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_43 <= line_shift_15_r_42; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_44 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_44 <= line_shift_15_r_43; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_45 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_45 <= line_shift_15_r_44; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_46 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_46 <= line_shift_15_r_45; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_47 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_47 <= line_shift_15_r_46; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_48 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_48 <= line_shift_15_r_47; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_49 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_49 <= line_shift_15_r_48; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_50 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_50 <= line_shift_15_r_49; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_51 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_51 <= line_shift_15_r_50; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_52 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_52 <= line_shift_15_r_51; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_53 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_53 <= line_shift_15_r_52; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_54 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_54 <= line_shift_15_r_53; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_55 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_55 <= line_shift_15_r_54; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_56 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_56 <= line_shift_15_r_55; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_57 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_57 <= line_shift_15_r_56; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_58 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_58 <= line_shift_15_r_57; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_59 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_59 <= line_shift_15_r_58; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_60 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_60 <= line_shift_15_r_59; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_61 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_61 <= line_shift_15_r_60; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_62 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_62 <= line_shift_15_r_61; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_63 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_63 <= line_shift_15_r_62; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_64 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_64 <= line_shift_15_r_63; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_65 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_65 <= line_shift_15_r_64; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_66 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_66 <= line_shift_15_r_65; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_67 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_67 <= line_shift_15_r_66; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_68 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_68 <= line_shift_15_r_67; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_69 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_69 <= line_shift_15_r_68; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_70 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_70 <= line_shift_15_r_69; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_71 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_71 <= line_shift_15_r_70; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_72 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_72 <= line_shift_15_r_71; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_73 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_73 <= line_shift_15_r_72; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_74 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_74 <= line_shift_15_r_73; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_75 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_75 <= line_shift_15_r_74; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_76 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_76 <= line_shift_15_r_75; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_77 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_77 <= line_shift_15_r_76; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_78 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_78 <= line_shift_15_r_77; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_79 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_79 <= line_shift_15_r_78; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_80 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_80 <= line_shift_15_r_79; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_81 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_81 <= line_shift_15_r_80; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_82 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_82 <= line_shift_15_r_81; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_83 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_83 <= line_shift_15_r_82; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_84 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_84 <= line_shift_15_r_83; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_85 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_85 <= line_shift_15_r_84; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_86 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_86 <= line_shift_15_r_85; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_87 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_87 <= line_shift_15_r_86; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_88 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_88 <= line_shift_15_r_87; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_89 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_89 <= line_shift_15_r_88; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_90 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_90 <= line_shift_15_r_89; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_91 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_91 <= line_shift_15_r_90; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_92 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_92 <= line_shift_15_r_91; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_93 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_93 <= line_shift_15_r_92; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_94 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_94 <= line_shift_15_r_93; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_95 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_95 <= line_shift_15_r_94; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_96 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_96 <= line_shift_15_r_95; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_97 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_97 <= line_shift_15_r_96; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_98 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_98 <= line_shift_15_r_97; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_99 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_99 <= line_shift_15_r_98; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_100 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_100 <= line_shift_15_r_99; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_101 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_101 <= line_shift_15_r_100; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_102 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_102 <= line_shift_15_r_101; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_103 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_103 <= line_shift_15_r_102; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_104 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_104 <= line_shift_15_r_103; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_105 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_105 <= line_shift_15_r_104; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_106 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_106 <= line_shift_15_r_105; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_107 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_107 <= line_shift_15_r_106; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_108 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_108 <= line_shift_15_r_107; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_109 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_109 <= line_shift_15_r_108; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_110 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_110 <= line_shift_15_r_109; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_111 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_111 <= line_shift_15_r_110; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_112 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_112 <= line_shift_15_r_111; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_113 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_113 <= line_shift_15_r_112; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_114 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_114 <= line_shift_15_r_113; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_115 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_115 <= line_shift_15_r_114; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_116 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_116 <= line_shift_15_r_115; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_117 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_117 <= line_shift_15_r_116; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_118 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_118 <= line_shift_15_r_117; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_119 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_119 <= line_shift_15_r_118; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_120 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_120 <= line_shift_15_r_119; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_121 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_121 <= line_shift_15_r_120; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_122 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_122 <= line_shift_15_r_121; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_123 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_123 <= line_shift_15_r_122; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_124 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_124 <= line_shift_15_r_123; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_125 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_125 <= line_shift_15_r_124; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_126 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_126 <= line_shift_15_r_125; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_127 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_127 <= line_shift_15_r_126; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_128 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_128 <= line_shift_15_r_127; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_129 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_129 <= line_shift_15_r_128; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_130 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_130 <= line_shift_15_r_129; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_131 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_131 <= line_shift_15_r_130; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_132 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_132 <= line_shift_15_r_131; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_133 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_133 <= line_shift_15_r_132; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_134 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_134 <= line_shift_15_r_133; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_135 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_135 <= line_shift_15_r_134; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_136 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_136 <= line_shift_15_r_135; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_137 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_137 <= line_shift_15_r_136; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_138 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_138 <= line_shift_15_r_137; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_139 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_139 <= line_shift_15_r_138; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_140 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_140 <= line_shift_15_r_139; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_141 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_141 <= line_shift_15_r_140; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_142 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_142 <= line_shift_15_r_141; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_143 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_143 <= line_shift_15_r_142; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_144 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_144 <= line_shift_15_r_143; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_145 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_145 <= line_shift_15_r_144; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_146 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_146 <= line_shift_15_r_145; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_147 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_147 <= line_shift_15_r_146; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_148 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_148 <= line_shift_15_r_147; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_149 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_149 <= line_shift_15_r_148; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_150 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_150 <= line_shift_15_r_149; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_151 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_151 <= line_shift_15_r_150; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_152 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_152 <= line_shift_15_r_151; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_153 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_153 <= line_shift_15_r_152; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_154 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_154 <= line_shift_15_r_153; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_155 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_155 <= line_shift_15_r_154; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_156 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_156 <= line_shift_15_r_155; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_157 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_157 <= line_shift_15_r_156; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15_r_158 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15_r_158 <= line_shift_15_r_157; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_line_extend_en) begin // @[Reg.scala 36:18]
      line_shift_15 <= line_shift_15_r_158; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_temp0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  reg_temp1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  reg_temp2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  line_shift_1_r = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  line_shift_1_r_1 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  line_shift_1_r_2 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  line_shift_1_r_3 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  line_shift_1_r_4 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  line_shift_1_r_5 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  line_shift_1_r_6 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  line_shift_1_r_7 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  line_shift_1_r_8 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  line_shift_1_r_9 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  line_shift_1_r_10 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  line_shift_1_r_11 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  line_shift_1_r_12 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  line_shift_1_r_13 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  line_shift_1_r_14 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  line_shift_1_r_15 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  line_shift_1_r_16 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  line_shift_1_r_17 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  line_shift_1_r_18 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  line_shift_1 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  line_shift_2_r = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  line_shift_2_r_1 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  line_shift_2_r_2 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  line_shift_2_r_3 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  line_shift_2_r_4 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  line_shift_2_r_5 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  line_shift_2_r_6 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  line_shift_2_r_7 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  line_shift_2_r_8 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  line_shift_2_r_9 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  line_shift_2_r_10 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  line_shift_2_r_11 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  line_shift_2_r_12 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  line_shift_2_r_13 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  line_shift_2_r_14 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  line_shift_2_r_15 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  line_shift_2_r_16 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  line_shift_2_r_17 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  line_shift_2_r_18 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  line_shift_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  line_shift_3_r = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  line_shift_3_r_1 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  line_shift_3_r_2 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  line_shift_3_r_3 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  line_shift_3_r_4 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  line_shift_3_r_5 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  line_shift_3_r_6 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  line_shift_3_r_7 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  line_shift_3_r_8 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  line_shift_3_r_9 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  line_shift_3_r_10 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  line_shift_3_r_11 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  line_shift_3_r_12 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  line_shift_3_r_13 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  line_shift_3_r_14 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  line_shift_3_r_15 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  line_shift_3_r_16 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  line_shift_3_r_17 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  line_shift_3_r_18 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  line_shift_3_r_19 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  line_shift_3_r_20 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  line_shift_3_r_21 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  line_shift_3_r_22 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  line_shift_3_r_23 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  line_shift_3_r_24 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  line_shift_3_r_25 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  line_shift_3_r_26 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  line_shift_3_r_27 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  line_shift_3_r_28 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  line_shift_3_r_29 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  line_shift_3_r_30 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  line_shift_3_r_31 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  line_shift_3_r_32 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  line_shift_3_r_33 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  line_shift_3_r_34 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  line_shift_3_r_35 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  line_shift_3_r_36 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  line_shift_3_r_37 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  line_shift_3_r_38 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  line_shift_3 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  line_shift_4_r = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  line_shift_4_r_1 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  line_shift_4_r_2 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  line_shift_4_r_3 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  line_shift_4_r_4 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  line_shift_4_r_5 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  line_shift_4_r_6 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  line_shift_4_r_7 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  line_shift_4_r_8 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  line_shift_4_r_9 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  line_shift_4_r_10 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  line_shift_4_r_11 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  line_shift_4_r_12 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  line_shift_4_r_13 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  line_shift_4_r_14 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  line_shift_4_r_15 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  line_shift_4_r_16 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  line_shift_4_r_17 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  line_shift_4_r_18 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  line_shift_4_r_19 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  line_shift_4_r_20 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  line_shift_4_r_21 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  line_shift_4_r_22 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  line_shift_4_r_23 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  line_shift_4_r_24 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  line_shift_4_r_25 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  line_shift_4_r_26 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  line_shift_4_r_27 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  line_shift_4_r_28 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  line_shift_4_r_29 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  line_shift_4_r_30 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  line_shift_4_r_31 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  line_shift_4_r_32 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  line_shift_4_r_33 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  line_shift_4_r_34 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  line_shift_4_r_35 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  line_shift_4_r_36 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  line_shift_4_r_37 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  line_shift_4_r_38 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  line_shift_4_r_39 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  line_shift_4_r_40 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  line_shift_4_r_41 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  line_shift_4_r_42 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  line_shift_4_r_43 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  line_shift_4_r_44 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  line_shift_4_r_45 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  line_shift_4_r_46 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  line_shift_4_r_47 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  line_shift_4_r_48 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  line_shift_4_r_49 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  line_shift_4_r_50 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  line_shift_4_r_51 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  line_shift_4_r_52 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  line_shift_4_r_53 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  line_shift_4_r_54 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  line_shift_4_r_55 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  line_shift_4_r_56 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  line_shift_4_r_57 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  line_shift_4_r_58 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  line_shift_4_r_59 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  line_shift_4_r_60 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  line_shift_4_r_61 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  line_shift_4_r_62 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  line_shift_4_r_63 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  line_shift_4_r_64 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  line_shift_4_r_65 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  line_shift_4_r_66 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  line_shift_4_r_67 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  line_shift_4_r_68 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  line_shift_4_r_69 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  line_shift_4_r_70 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  line_shift_4_r_71 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  line_shift_4_r_72 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  line_shift_4_r_73 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  line_shift_4_r_74 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  line_shift_4_r_75 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  line_shift_4_r_76 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  line_shift_4_r_77 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  line_shift_4_r_78 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  line_shift_4 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  line_shift_5_r = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  line_shift_5_r_1 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  line_shift_5_r_2 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  line_shift_5_r_3 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  line_shift_5_r_4 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  line_shift_5_r_5 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  line_shift_5_r_6 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  line_shift_5_r_7 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  line_shift_5_r_8 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  line_shift_5_r_9 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  line_shift_5_r_10 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  line_shift_5_r_11 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  line_shift_5_r_12 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  line_shift_5_r_13 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  line_shift_5_r_14 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  line_shift_5_r_15 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  line_shift_5_r_16 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  line_shift_5_r_17 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  line_shift_5_r_18 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  line_shift_5_r_19 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  line_shift_5_r_20 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  line_shift_5_r_21 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  line_shift_5_r_22 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  line_shift_5_r_23 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  line_shift_5_r_24 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  line_shift_5_r_25 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  line_shift_5_r_26 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  line_shift_5_r_27 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  line_shift_5_r_28 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  line_shift_5_r_29 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  line_shift_5_r_30 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  line_shift_5_r_31 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  line_shift_5_r_32 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  line_shift_5_r_33 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  line_shift_5_r_34 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  line_shift_5_r_35 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  line_shift_5_r_36 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  line_shift_5_r_37 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  line_shift_5_r_38 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  line_shift_5_r_39 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  line_shift_5_r_40 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  line_shift_5_r_41 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  line_shift_5_r_42 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  line_shift_5_r_43 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  line_shift_5_r_44 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  line_shift_5_r_45 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  line_shift_5_r_46 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  line_shift_5_r_47 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  line_shift_5_r_48 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  line_shift_5_r_49 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  line_shift_5_r_50 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  line_shift_5_r_51 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  line_shift_5_r_52 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  line_shift_5_r_53 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  line_shift_5_r_54 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  line_shift_5_r_55 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  line_shift_5_r_56 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  line_shift_5_r_57 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  line_shift_5_r_58 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  line_shift_5_r_59 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  line_shift_5_r_60 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  line_shift_5_r_61 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  line_shift_5_r_62 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  line_shift_5_r_63 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  line_shift_5_r_64 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  line_shift_5_r_65 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  line_shift_5_r_66 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  line_shift_5_r_67 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  line_shift_5_r_68 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  line_shift_5_r_69 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  line_shift_5_r_70 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  line_shift_5_r_71 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  line_shift_5_r_72 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  line_shift_5_r_73 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  line_shift_5_r_74 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  line_shift_5_r_75 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  line_shift_5_r_76 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  line_shift_5_r_77 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  line_shift_5_r_78 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  line_shift_5_r_79 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  line_shift_5_r_80 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  line_shift_5_r_81 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  line_shift_5_r_82 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  line_shift_5_r_83 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  line_shift_5_r_84 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  line_shift_5_r_85 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  line_shift_5_r_86 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  line_shift_5_r_87 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  line_shift_5_r_88 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  line_shift_5_r_89 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  line_shift_5_r_90 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  line_shift_5_r_91 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  line_shift_5_r_92 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  line_shift_5_r_93 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  line_shift_5_r_94 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  line_shift_5_r_95 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  line_shift_5_r_96 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  line_shift_5_r_97 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  line_shift_5_r_98 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  line_shift_5_r_99 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  line_shift_5_r_100 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  line_shift_5_r_101 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  line_shift_5_r_102 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  line_shift_5_r_103 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  line_shift_5_r_104 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  line_shift_5_r_105 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  line_shift_5_r_106 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  line_shift_5_r_107 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  line_shift_5_r_108 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  line_shift_5_r_109 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  line_shift_5_r_110 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  line_shift_5_r_111 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  line_shift_5_r_112 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  line_shift_5_r_113 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  line_shift_5_r_114 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  line_shift_5_r_115 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  line_shift_5_r_116 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  line_shift_5_r_117 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  line_shift_5_r_118 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  line_shift_5_r_119 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  line_shift_5_r_120 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  line_shift_5_r_121 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  line_shift_5_r_122 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  line_shift_5_r_123 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  line_shift_5_r_124 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  line_shift_5_r_125 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  line_shift_5_r_126 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  line_shift_5_r_127 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  line_shift_5_r_128 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  line_shift_5_r_129 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  line_shift_5_r_130 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  line_shift_5_r_131 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  line_shift_5_r_132 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  line_shift_5_r_133 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  line_shift_5_r_134 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  line_shift_5_r_135 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  line_shift_5_r_136 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  line_shift_5_r_137 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  line_shift_5_r_138 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  line_shift_5_r_139 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  line_shift_5_r_140 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  line_shift_5_r_141 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  line_shift_5_r_142 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  line_shift_5_r_143 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  line_shift_5_r_144 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  line_shift_5_r_145 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  line_shift_5_r_146 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  line_shift_5_r_147 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  line_shift_5_r_148 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  line_shift_5_r_149 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  line_shift_5_r_150 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  line_shift_5_r_151 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  line_shift_5_r_152 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  line_shift_5_r_153 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  line_shift_5_r_154 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  line_shift_5_r_155 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  line_shift_5_r_156 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  line_shift_5_r_157 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  line_shift_5_r_158 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  line_shift_5 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  line_shift_11_r = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  line_shift_11_r_1 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  line_shift_11_r_2 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  line_shift_11_r_3 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  line_shift_11_r_4 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  line_shift_11_r_5 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  line_shift_11_r_6 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  line_shift_11_r_7 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  line_shift_11_r_8 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  line_shift_11_r_9 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  line_shift_11_r_10 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  line_shift_11_r_11 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  line_shift_11_r_12 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  line_shift_11_r_13 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  line_shift_11_r_14 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  line_shift_11_r_15 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  line_shift_11_r_16 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  line_shift_11_r_17 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  line_shift_11_r_18 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  line_shift_11 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  line_shift_12_r = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  line_shift_12_r_1 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  line_shift_12_r_2 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  line_shift_12_r_3 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  line_shift_12_r_4 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  line_shift_12_r_5 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  line_shift_12_r_6 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  line_shift_12_r_7 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  line_shift_12_r_8 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  line_shift_12_r_9 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  line_shift_12_r_10 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  line_shift_12_r_11 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  line_shift_12_r_12 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  line_shift_12_r_13 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  line_shift_12_r_14 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  line_shift_12_r_15 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  line_shift_12_r_16 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  line_shift_12_r_17 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  line_shift_12_r_18 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  line_shift_12 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  line_shift_13_r = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  line_shift_13_r_1 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  line_shift_13_r_2 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  line_shift_13_r_3 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  line_shift_13_r_4 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  line_shift_13_r_5 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  line_shift_13_r_6 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  line_shift_13_r_7 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  line_shift_13_r_8 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  line_shift_13_r_9 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  line_shift_13_r_10 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  line_shift_13_r_11 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  line_shift_13_r_12 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  line_shift_13_r_13 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  line_shift_13_r_14 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  line_shift_13_r_15 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  line_shift_13_r_16 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  line_shift_13_r_17 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  line_shift_13_r_18 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  line_shift_13_r_19 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  line_shift_13_r_20 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  line_shift_13_r_21 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  line_shift_13_r_22 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  line_shift_13_r_23 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  line_shift_13_r_24 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  line_shift_13_r_25 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  line_shift_13_r_26 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  line_shift_13_r_27 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  line_shift_13_r_28 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  line_shift_13_r_29 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  line_shift_13_r_30 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  line_shift_13_r_31 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  line_shift_13_r_32 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  line_shift_13_r_33 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  line_shift_13_r_34 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  line_shift_13_r_35 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  line_shift_13_r_36 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  line_shift_13_r_37 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  line_shift_13_r_38 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  line_shift_13 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  line_shift_14_r = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  line_shift_14_r_1 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  line_shift_14_r_2 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  line_shift_14_r_3 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  line_shift_14_r_4 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  line_shift_14_r_5 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  line_shift_14_r_6 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  line_shift_14_r_7 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  line_shift_14_r_8 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  line_shift_14_r_9 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  line_shift_14_r_10 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  line_shift_14_r_11 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  line_shift_14_r_12 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  line_shift_14_r_13 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  line_shift_14_r_14 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  line_shift_14_r_15 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  line_shift_14_r_16 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  line_shift_14_r_17 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  line_shift_14_r_18 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  line_shift_14_r_19 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  line_shift_14_r_20 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  line_shift_14_r_21 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  line_shift_14_r_22 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  line_shift_14_r_23 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  line_shift_14_r_24 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  line_shift_14_r_25 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  line_shift_14_r_26 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  line_shift_14_r_27 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  line_shift_14_r_28 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  line_shift_14_r_29 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  line_shift_14_r_30 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  line_shift_14_r_31 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  line_shift_14_r_32 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  line_shift_14_r_33 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  line_shift_14_r_34 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  line_shift_14_r_35 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  line_shift_14_r_36 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  line_shift_14_r_37 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  line_shift_14_r_38 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  line_shift_14_r_39 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  line_shift_14_r_40 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  line_shift_14_r_41 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  line_shift_14_r_42 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  line_shift_14_r_43 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  line_shift_14_r_44 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  line_shift_14_r_45 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  line_shift_14_r_46 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  line_shift_14_r_47 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  line_shift_14_r_48 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  line_shift_14_r_49 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  line_shift_14_r_50 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  line_shift_14_r_51 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  line_shift_14_r_52 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  line_shift_14_r_53 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  line_shift_14_r_54 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  line_shift_14_r_55 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  line_shift_14_r_56 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  line_shift_14_r_57 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  line_shift_14_r_58 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  line_shift_14_r_59 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  line_shift_14_r_60 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  line_shift_14_r_61 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  line_shift_14_r_62 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  line_shift_14_r_63 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  line_shift_14_r_64 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  line_shift_14_r_65 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  line_shift_14_r_66 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  line_shift_14_r_67 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  line_shift_14_r_68 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  line_shift_14_r_69 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  line_shift_14_r_70 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  line_shift_14_r_71 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  line_shift_14_r_72 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  line_shift_14_r_73 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  line_shift_14_r_74 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  line_shift_14_r_75 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  line_shift_14_r_76 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  line_shift_14_r_77 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  line_shift_14_r_78 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  line_shift_14 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  line_shift_15_r = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  line_shift_15_r_1 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  line_shift_15_r_2 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  line_shift_15_r_3 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  line_shift_15_r_4 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  line_shift_15_r_5 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  line_shift_15_r_6 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  line_shift_15_r_7 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  line_shift_15_r_8 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  line_shift_15_r_9 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  line_shift_15_r_10 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  line_shift_15_r_11 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  line_shift_15_r_12 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  line_shift_15_r_13 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  line_shift_15_r_14 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  line_shift_15_r_15 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  line_shift_15_r_16 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  line_shift_15_r_17 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  line_shift_15_r_18 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  line_shift_15_r_19 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  line_shift_15_r_20 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  line_shift_15_r_21 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  line_shift_15_r_22 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  line_shift_15_r_23 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  line_shift_15_r_24 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  line_shift_15_r_25 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  line_shift_15_r_26 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  line_shift_15_r_27 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  line_shift_15_r_28 = _RAND_511[7:0];
  _RAND_512 = {1{`RANDOM}};
  line_shift_15_r_29 = _RAND_512[7:0];
  _RAND_513 = {1{`RANDOM}};
  line_shift_15_r_30 = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  line_shift_15_r_31 = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  line_shift_15_r_32 = _RAND_515[7:0];
  _RAND_516 = {1{`RANDOM}};
  line_shift_15_r_33 = _RAND_516[7:0];
  _RAND_517 = {1{`RANDOM}};
  line_shift_15_r_34 = _RAND_517[7:0];
  _RAND_518 = {1{`RANDOM}};
  line_shift_15_r_35 = _RAND_518[7:0];
  _RAND_519 = {1{`RANDOM}};
  line_shift_15_r_36 = _RAND_519[7:0];
  _RAND_520 = {1{`RANDOM}};
  line_shift_15_r_37 = _RAND_520[7:0];
  _RAND_521 = {1{`RANDOM}};
  line_shift_15_r_38 = _RAND_521[7:0];
  _RAND_522 = {1{`RANDOM}};
  line_shift_15_r_39 = _RAND_522[7:0];
  _RAND_523 = {1{`RANDOM}};
  line_shift_15_r_40 = _RAND_523[7:0];
  _RAND_524 = {1{`RANDOM}};
  line_shift_15_r_41 = _RAND_524[7:0];
  _RAND_525 = {1{`RANDOM}};
  line_shift_15_r_42 = _RAND_525[7:0];
  _RAND_526 = {1{`RANDOM}};
  line_shift_15_r_43 = _RAND_526[7:0];
  _RAND_527 = {1{`RANDOM}};
  line_shift_15_r_44 = _RAND_527[7:0];
  _RAND_528 = {1{`RANDOM}};
  line_shift_15_r_45 = _RAND_528[7:0];
  _RAND_529 = {1{`RANDOM}};
  line_shift_15_r_46 = _RAND_529[7:0];
  _RAND_530 = {1{`RANDOM}};
  line_shift_15_r_47 = _RAND_530[7:0];
  _RAND_531 = {1{`RANDOM}};
  line_shift_15_r_48 = _RAND_531[7:0];
  _RAND_532 = {1{`RANDOM}};
  line_shift_15_r_49 = _RAND_532[7:0];
  _RAND_533 = {1{`RANDOM}};
  line_shift_15_r_50 = _RAND_533[7:0];
  _RAND_534 = {1{`RANDOM}};
  line_shift_15_r_51 = _RAND_534[7:0];
  _RAND_535 = {1{`RANDOM}};
  line_shift_15_r_52 = _RAND_535[7:0];
  _RAND_536 = {1{`RANDOM}};
  line_shift_15_r_53 = _RAND_536[7:0];
  _RAND_537 = {1{`RANDOM}};
  line_shift_15_r_54 = _RAND_537[7:0];
  _RAND_538 = {1{`RANDOM}};
  line_shift_15_r_55 = _RAND_538[7:0];
  _RAND_539 = {1{`RANDOM}};
  line_shift_15_r_56 = _RAND_539[7:0];
  _RAND_540 = {1{`RANDOM}};
  line_shift_15_r_57 = _RAND_540[7:0];
  _RAND_541 = {1{`RANDOM}};
  line_shift_15_r_58 = _RAND_541[7:0];
  _RAND_542 = {1{`RANDOM}};
  line_shift_15_r_59 = _RAND_542[7:0];
  _RAND_543 = {1{`RANDOM}};
  line_shift_15_r_60 = _RAND_543[7:0];
  _RAND_544 = {1{`RANDOM}};
  line_shift_15_r_61 = _RAND_544[7:0];
  _RAND_545 = {1{`RANDOM}};
  line_shift_15_r_62 = _RAND_545[7:0];
  _RAND_546 = {1{`RANDOM}};
  line_shift_15_r_63 = _RAND_546[7:0];
  _RAND_547 = {1{`RANDOM}};
  line_shift_15_r_64 = _RAND_547[7:0];
  _RAND_548 = {1{`RANDOM}};
  line_shift_15_r_65 = _RAND_548[7:0];
  _RAND_549 = {1{`RANDOM}};
  line_shift_15_r_66 = _RAND_549[7:0];
  _RAND_550 = {1{`RANDOM}};
  line_shift_15_r_67 = _RAND_550[7:0];
  _RAND_551 = {1{`RANDOM}};
  line_shift_15_r_68 = _RAND_551[7:0];
  _RAND_552 = {1{`RANDOM}};
  line_shift_15_r_69 = _RAND_552[7:0];
  _RAND_553 = {1{`RANDOM}};
  line_shift_15_r_70 = _RAND_553[7:0];
  _RAND_554 = {1{`RANDOM}};
  line_shift_15_r_71 = _RAND_554[7:0];
  _RAND_555 = {1{`RANDOM}};
  line_shift_15_r_72 = _RAND_555[7:0];
  _RAND_556 = {1{`RANDOM}};
  line_shift_15_r_73 = _RAND_556[7:0];
  _RAND_557 = {1{`RANDOM}};
  line_shift_15_r_74 = _RAND_557[7:0];
  _RAND_558 = {1{`RANDOM}};
  line_shift_15_r_75 = _RAND_558[7:0];
  _RAND_559 = {1{`RANDOM}};
  line_shift_15_r_76 = _RAND_559[7:0];
  _RAND_560 = {1{`RANDOM}};
  line_shift_15_r_77 = _RAND_560[7:0];
  _RAND_561 = {1{`RANDOM}};
  line_shift_15_r_78 = _RAND_561[7:0];
  _RAND_562 = {1{`RANDOM}};
  line_shift_15_r_79 = _RAND_562[7:0];
  _RAND_563 = {1{`RANDOM}};
  line_shift_15_r_80 = _RAND_563[7:0];
  _RAND_564 = {1{`RANDOM}};
  line_shift_15_r_81 = _RAND_564[7:0];
  _RAND_565 = {1{`RANDOM}};
  line_shift_15_r_82 = _RAND_565[7:0];
  _RAND_566 = {1{`RANDOM}};
  line_shift_15_r_83 = _RAND_566[7:0];
  _RAND_567 = {1{`RANDOM}};
  line_shift_15_r_84 = _RAND_567[7:0];
  _RAND_568 = {1{`RANDOM}};
  line_shift_15_r_85 = _RAND_568[7:0];
  _RAND_569 = {1{`RANDOM}};
  line_shift_15_r_86 = _RAND_569[7:0];
  _RAND_570 = {1{`RANDOM}};
  line_shift_15_r_87 = _RAND_570[7:0];
  _RAND_571 = {1{`RANDOM}};
  line_shift_15_r_88 = _RAND_571[7:0];
  _RAND_572 = {1{`RANDOM}};
  line_shift_15_r_89 = _RAND_572[7:0];
  _RAND_573 = {1{`RANDOM}};
  line_shift_15_r_90 = _RAND_573[7:0];
  _RAND_574 = {1{`RANDOM}};
  line_shift_15_r_91 = _RAND_574[7:0];
  _RAND_575 = {1{`RANDOM}};
  line_shift_15_r_92 = _RAND_575[7:0];
  _RAND_576 = {1{`RANDOM}};
  line_shift_15_r_93 = _RAND_576[7:0];
  _RAND_577 = {1{`RANDOM}};
  line_shift_15_r_94 = _RAND_577[7:0];
  _RAND_578 = {1{`RANDOM}};
  line_shift_15_r_95 = _RAND_578[7:0];
  _RAND_579 = {1{`RANDOM}};
  line_shift_15_r_96 = _RAND_579[7:0];
  _RAND_580 = {1{`RANDOM}};
  line_shift_15_r_97 = _RAND_580[7:0];
  _RAND_581 = {1{`RANDOM}};
  line_shift_15_r_98 = _RAND_581[7:0];
  _RAND_582 = {1{`RANDOM}};
  line_shift_15_r_99 = _RAND_582[7:0];
  _RAND_583 = {1{`RANDOM}};
  line_shift_15_r_100 = _RAND_583[7:0];
  _RAND_584 = {1{`RANDOM}};
  line_shift_15_r_101 = _RAND_584[7:0];
  _RAND_585 = {1{`RANDOM}};
  line_shift_15_r_102 = _RAND_585[7:0];
  _RAND_586 = {1{`RANDOM}};
  line_shift_15_r_103 = _RAND_586[7:0];
  _RAND_587 = {1{`RANDOM}};
  line_shift_15_r_104 = _RAND_587[7:0];
  _RAND_588 = {1{`RANDOM}};
  line_shift_15_r_105 = _RAND_588[7:0];
  _RAND_589 = {1{`RANDOM}};
  line_shift_15_r_106 = _RAND_589[7:0];
  _RAND_590 = {1{`RANDOM}};
  line_shift_15_r_107 = _RAND_590[7:0];
  _RAND_591 = {1{`RANDOM}};
  line_shift_15_r_108 = _RAND_591[7:0];
  _RAND_592 = {1{`RANDOM}};
  line_shift_15_r_109 = _RAND_592[7:0];
  _RAND_593 = {1{`RANDOM}};
  line_shift_15_r_110 = _RAND_593[7:0];
  _RAND_594 = {1{`RANDOM}};
  line_shift_15_r_111 = _RAND_594[7:0];
  _RAND_595 = {1{`RANDOM}};
  line_shift_15_r_112 = _RAND_595[7:0];
  _RAND_596 = {1{`RANDOM}};
  line_shift_15_r_113 = _RAND_596[7:0];
  _RAND_597 = {1{`RANDOM}};
  line_shift_15_r_114 = _RAND_597[7:0];
  _RAND_598 = {1{`RANDOM}};
  line_shift_15_r_115 = _RAND_598[7:0];
  _RAND_599 = {1{`RANDOM}};
  line_shift_15_r_116 = _RAND_599[7:0];
  _RAND_600 = {1{`RANDOM}};
  line_shift_15_r_117 = _RAND_600[7:0];
  _RAND_601 = {1{`RANDOM}};
  line_shift_15_r_118 = _RAND_601[7:0];
  _RAND_602 = {1{`RANDOM}};
  line_shift_15_r_119 = _RAND_602[7:0];
  _RAND_603 = {1{`RANDOM}};
  line_shift_15_r_120 = _RAND_603[7:0];
  _RAND_604 = {1{`RANDOM}};
  line_shift_15_r_121 = _RAND_604[7:0];
  _RAND_605 = {1{`RANDOM}};
  line_shift_15_r_122 = _RAND_605[7:0];
  _RAND_606 = {1{`RANDOM}};
  line_shift_15_r_123 = _RAND_606[7:0];
  _RAND_607 = {1{`RANDOM}};
  line_shift_15_r_124 = _RAND_607[7:0];
  _RAND_608 = {1{`RANDOM}};
  line_shift_15_r_125 = _RAND_608[7:0];
  _RAND_609 = {1{`RANDOM}};
  line_shift_15_r_126 = _RAND_609[7:0];
  _RAND_610 = {1{`RANDOM}};
  line_shift_15_r_127 = _RAND_610[7:0];
  _RAND_611 = {1{`RANDOM}};
  line_shift_15_r_128 = _RAND_611[7:0];
  _RAND_612 = {1{`RANDOM}};
  line_shift_15_r_129 = _RAND_612[7:0];
  _RAND_613 = {1{`RANDOM}};
  line_shift_15_r_130 = _RAND_613[7:0];
  _RAND_614 = {1{`RANDOM}};
  line_shift_15_r_131 = _RAND_614[7:0];
  _RAND_615 = {1{`RANDOM}};
  line_shift_15_r_132 = _RAND_615[7:0];
  _RAND_616 = {1{`RANDOM}};
  line_shift_15_r_133 = _RAND_616[7:0];
  _RAND_617 = {1{`RANDOM}};
  line_shift_15_r_134 = _RAND_617[7:0];
  _RAND_618 = {1{`RANDOM}};
  line_shift_15_r_135 = _RAND_618[7:0];
  _RAND_619 = {1{`RANDOM}};
  line_shift_15_r_136 = _RAND_619[7:0];
  _RAND_620 = {1{`RANDOM}};
  line_shift_15_r_137 = _RAND_620[7:0];
  _RAND_621 = {1{`RANDOM}};
  line_shift_15_r_138 = _RAND_621[7:0];
  _RAND_622 = {1{`RANDOM}};
  line_shift_15_r_139 = _RAND_622[7:0];
  _RAND_623 = {1{`RANDOM}};
  line_shift_15_r_140 = _RAND_623[7:0];
  _RAND_624 = {1{`RANDOM}};
  line_shift_15_r_141 = _RAND_624[7:0];
  _RAND_625 = {1{`RANDOM}};
  line_shift_15_r_142 = _RAND_625[7:0];
  _RAND_626 = {1{`RANDOM}};
  line_shift_15_r_143 = _RAND_626[7:0];
  _RAND_627 = {1{`RANDOM}};
  line_shift_15_r_144 = _RAND_627[7:0];
  _RAND_628 = {1{`RANDOM}};
  line_shift_15_r_145 = _RAND_628[7:0];
  _RAND_629 = {1{`RANDOM}};
  line_shift_15_r_146 = _RAND_629[7:0];
  _RAND_630 = {1{`RANDOM}};
  line_shift_15_r_147 = _RAND_630[7:0];
  _RAND_631 = {1{`RANDOM}};
  line_shift_15_r_148 = _RAND_631[7:0];
  _RAND_632 = {1{`RANDOM}};
  line_shift_15_r_149 = _RAND_632[7:0];
  _RAND_633 = {1{`RANDOM}};
  line_shift_15_r_150 = _RAND_633[7:0];
  _RAND_634 = {1{`RANDOM}};
  line_shift_15_r_151 = _RAND_634[7:0];
  _RAND_635 = {1{`RANDOM}};
  line_shift_15_r_152 = _RAND_635[7:0];
  _RAND_636 = {1{`RANDOM}};
  line_shift_15_r_153 = _RAND_636[7:0];
  _RAND_637 = {1{`RANDOM}};
  line_shift_15_r_154 = _RAND_637[7:0];
  _RAND_638 = {1{`RANDOM}};
  line_shift_15_r_155 = _RAND_638[7:0];
  _RAND_639 = {1{`RANDOM}};
  line_shift_15_r_156 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  line_shift_15_r_157 = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  line_shift_15_r_158 = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  line_shift_15 = _RAND_642[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module line_buffer_unit_extend(
  input         clock,
  input         reset,
  input  [2:0]  io_sel,
  input         io_s_mod,
  input  [31:0] io_line_i_data,
  output [7:0]  io_line_o_data_0,
  output [7:0]  io_line_o_data_1,
  output [7:0]  io_line_o_data_2,
  output [7:0]  io_line_o_data_3,
  output [7:0]  io_line_o_data_4,
  output [7:0]  io_line_o_data_5,
  output [7:0]  io_line_o_data_6,
  output [7:0]  io_line_o_data_7,
  output [7:0]  io_line_o_data_8
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  line_0_clock; // @[LineBuffer.scala 159:34]
  wire  line_0_reset; // @[LineBuffer.scala 159:34]
  wire [15:0] line_0_io_i; // @[LineBuffer.scala 159:34]
  wire [15:0] line_0_io_o; // @[LineBuffer.scala 159:34]
  wire  line_0_io_s_mod; // @[LineBuffer.scala 159:34]
  wire  line_0_io_line_extend_en; // @[LineBuffer.scala 159:34]
  wire [2:0] line_0_io_sel; // @[LineBuffer.scala 159:34]
  wire  line_1_clock; // @[LineBuffer.scala 159:34]
  wire  line_1_reset; // @[LineBuffer.scala 159:34]
  wire [15:0] line_1_io_i; // @[LineBuffer.scala 159:34]
  wire [15:0] line_1_io_o; // @[LineBuffer.scala 159:34]
  wire  line_1_io_s_mod; // @[LineBuffer.scala 159:34]
  wire  line_1_io_line_extend_en; // @[LineBuffer.scala 159:34]
  wire [2:0] line_1_io_sel; // @[LineBuffer.scala 159:34]
  reg [7:0] win_0; // @[LineBuffer.scala 174:34]
  reg [7:0] win_1; // @[LineBuffer.scala 174:34]
  reg [7:0] win_2; // @[LineBuffer.scala 174:34]
  reg [7:0] win_3; // @[LineBuffer.scala 174:34]
  reg [7:0] win_4; // @[LineBuffer.scala 174:34]
  reg [7:0] win_5; // @[LineBuffer.scala 174:34]
  reg [7:0] win_6; // @[LineBuffer.scala 174:34]
  reg [7:0] win_7; // @[LineBuffer.scala 174:34]
  reg [7:0] win_8; // @[LineBuffer.scala 174:34]
  wire [15:0] line_out_0 = line_1_io_o; // @[LineBuffer.scala 169:24 170:17]
  wire [15:0] line_out_1 = line_0_io_o; // @[LineBuffer.scala 169:24 171:17]
  reg [7:0] temp_win_0; // @[LineBuffer.scala 187:39]
  reg [7:0] temp_win_1; // @[LineBuffer.scala 187:39]
  reg [7:0] temp_win_2; // @[LineBuffer.scala 187:39]
  linebuf_unit_extend line_0 ( // @[LineBuffer.scala 159:34]
    .clock(line_0_clock),
    .reset(line_0_reset),
    .io_i(line_0_io_i),
    .io_o(line_0_io_o),
    .io_s_mod(line_0_io_s_mod),
    .io_line_extend_en(line_0_io_line_extend_en),
    .io_sel(line_0_io_sel)
  );
  linebuf_unit_extend line_1 ( // @[LineBuffer.scala 159:34]
    .clock(line_1_clock),
    .reset(line_1_reset),
    .io_i(line_1_io_i),
    .io_o(line_1_io_o),
    .io_s_mod(line_1_io_s_mod),
    .io_line_extend_en(line_1_io_line_extend_en),
    .io_sel(line_1_io_sel)
  );
  assign io_line_o_data_0 = io_s_mod ? temp_win_0 : win_0; // @[LineBuffer.scala 192:29]
  assign io_line_o_data_1 = io_s_mod ? win_0 : win_1; // @[LineBuffer.scala 193:29]
  assign io_line_o_data_2 = io_s_mod ? win_1 : win_2; // @[LineBuffer.scala 194:29]
  assign io_line_o_data_3 = io_s_mod ? temp_win_1 : win_3; // @[LineBuffer.scala 195:29]
  assign io_line_o_data_4 = io_s_mod ? win_3 : win_4; // @[LineBuffer.scala 196:29]
  assign io_line_o_data_5 = io_s_mod ? win_4 : win_5; // @[LineBuffer.scala 197:29]
  assign io_line_o_data_6 = io_s_mod ? temp_win_2 : win_6; // @[LineBuffer.scala 198:29]
  assign io_line_o_data_7 = io_s_mod ? win_6 : win_7; // @[LineBuffer.scala 199:29]
  assign io_line_o_data_8 = io_s_mod ? win_7 : win_8; // @[LineBuffer.scala 200:29]
  assign line_0_clock = clock;
  assign line_0_reset = reset;
  assign line_0_io_i = io_s_mod ? io_line_i_data[31:16] : io_line_i_data[15:0]; // @[LineBuffer.scala 168:24]
  assign line_0_io_s_mod = io_s_mod; // @[LineBuffer.scala 162:26]
  assign line_0_io_line_extend_en = io_s_mod; // @[LineBuffer.scala 158:27]
  assign line_0_io_sel = io_sel; // @[LineBuffer.scala 161:24]
  assign line_1_clock = clock;
  assign line_1_reset = reset;
  assign line_1_io_i = io_s_mod ? io_line_i_data[15:0] : line_0_io_o; // @[LineBuffer.scala 167:24]
  assign line_1_io_s_mod = io_s_mod; // @[LineBuffer.scala 162:26]
  assign line_1_io_line_extend_en = io_s_mod; // @[LineBuffer.scala 158:27]
  assign line_1_io_sel = io_sel; // @[LineBuffer.scala 161:24]
  always @(posedge clock) begin
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_0 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 175:18]
      win_0 <= win_2;
    end else begin
      win_0 <= win_1;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_1 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 179:18]
      win_1 <= line_out_0[7:0];
    end else begin
      win_1 <= win_2;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_2 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 183:18]
      win_2 <= line_out_0[15:8];
    end else begin
      win_2 <= line_out_0[7:0];
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_3 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 176:18]
      win_3 <= win_5;
    end else begin
      win_3 <= win_4;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_4 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 180:18]
      win_4 <= line_out_1[7:0];
    end else begin
      win_4 <= win_5;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_5 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 184:18]
      win_5 <= line_out_1[15:8];
    end else begin
      win_5 <= line_out_1[7:0];
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_6 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 177:18]
      win_6 <= win_8;
    end else begin
      win_6 <= win_7;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_7 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 181:18]
      win_7 <= io_line_i_data[7:0];
    end else begin
      win_7 <= win_8;
    end
    if (reset) begin // @[LineBuffer.scala 174:34]
      win_8 <= 8'h0; // @[LineBuffer.scala 174:34]
    end else if (io_s_mod) begin // @[LineBuffer.scala 185:18]
      win_8 <= io_line_i_data[15:8];
    end else begin
      win_8 <= io_line_i_data[7:0];
    end
    if (reset) begin // @[LineBuffer.scala 187:39]
      temp_win_0 <= 8'h0; // @[LineBuffer.scala 187:39]
    end else begin
      temp_win_0 <= win_1; // @[LineBuffer.scala 188:17]
    end
    if (reset) begin // @[LineBuffer.scala 187:39]
      temp_win_1 <= 8'h0; // @[LineBuffer.scala 187:39]
    end else begin
      temp_win_1 <= win_4; // @[LineBuffer.scala 189:17]
    end
    if (reset) begin // @[LineBuffer.scala 187:39]
      temp_win_2 <= 8'h0; // @[LineBuffer.scala 187:39]
    end else begin
      temp_win_2 <= win_7; // @[LineBuffer.scala 190:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  win_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  win_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  win_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  win_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  win_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  win_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  win_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  win_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  win_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  temp_win_0 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  temp_win_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  temp_win_2 = _RAND_11[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LineBuffer_extend(
  input         clock,
  input         reset,
  input  [2:0]  io_sel,
  input         io_s_mod,
  input  [31:0] io_lineBuffer_i_data_0,
  input  [31:0] io_lineBuffer_i_data_1,
  input  [31:0] io_lineBuffer_i_data_2,
  input  [31:0] io_lineBuffer_i_data_3,
  input  [31:0] io_lineBuffer_i_data_4,
  input  [31:0] io_lineBuffer_i_data_5,
  input  [31:0] io_lineBuffer_i_data_6,
  input  [31:0] io_lineBuffer_i_data_7,
  output [7:0]  io_lineBuffer_o_data_0,
  output [7:0]  io_lineBuffer_o_data_1,
  output [7:0]  io_lineBuffer_o_data_2,
  output [7:0]  io_lineBuffer_o_data_3,
  output [7:0]  io_lineBuffer_o_data_4,
  output [7:0]  io_lineBuffer_o_data_5,
  output [7:0]  io_lineBuffer_o_data_6,
  output [7:0]  io_lineBuffer_o_data_7,
  output [7:0]  io_lineBuffer_o_data_8,
  output [7:0]  io_lineBuffer_o_data_9,
  output [7:0]  io_lineBuffer_o_data_10,
  output [7:0]  io_lineBuffer_o_data_11,
  output [7:0]  io_lineBuffer_o_data_12,
  output [7:0]  io_lineBuffer_o_data_13,
  output [7:0]  io_lineBuffer_o_data_14,
  output [7:0]  io_lineBuffer_o_data_15,
  output [7:0]  io_lineBuffer_o_data_16,
  output [7:0]  io_lineBuffer_o_data_17,
  output [7:0]  io_lineBuffer_o_data_18,
  output [7:0]  io_lineBuffer_o_data_19,
  output [7:0]  io_lineBuffer_o_data_20,
  output [7:0]  io_lineBuffer_o_data_21,
  output [7:0]  io_lineBuffer_o_data_22,
  output [7:0]  io_lineBuffer_o_data_23,
  output [7:0]  io_lineBuffer_o_data_24,
  output [7:0]  io_lineBuffer_o_data_25,
  output [7:0]  io_lineBuffer_o_data_26,
  output [7:0]  io_lineBuffer_o_data_27,
  output [7:0]  io_lineBuffer_o_data_28,
  output [7:0]  io_lineBuffer_o_data_29,
  output [7:0]  io_lineBuffer_o_data_30,
  output [7:0]  io_lineBuffer_o_data_31,
  output [7:0]  io_lineBuffer_o_data_32,
  output [7:0]  io_lineBuffer_o_data_33,
  output [7:0]  io_lineBuffer_o_data_34,
  output [7:0]  io_lineBuffer_o_data_35,
  output [7:0]  io_lineBuffer_o_data_36,
  output [7:0]  io_lineBuffer_o_data_37,
  output [7:0]  io_lineBuffer_o_data_38,
  output [7:0]  io_lineBuffer_o_data_39,
  output [7:0]  io_lineBuffer_o_data_40,
  output [7:0]  io_lineBuffer_o_data_41,
  output [7:0]  io_lineBuffer_o_data_42,
  output [7:0]  io_lineBuffer_o_data_43,
  output [7:0]  io_lineBuffer_o_data_44,
  output [7:0]  io_lineBuffer_o_data_45,
  output [7:0]  io_lineBuffer_o_data_46,
  output [7:0]  io_lineBuffer_o_data_47,
  output [7:0]  io_lineBuffer_o_data_48,
  output [7:0]  io_lineBuffer_o_data_49,
  output [7:0]  io_lineBuffer_o_data_50,
  output [7:0]  io_lineBuffer_o_data_51,
  output [7:0]  io_lineBuffer_o_data_52,
  output [7:0]  io_lineBuffer_o_data_53,
  output [7:0]  io_lineBuffer_o_data_54,
  output [7:0]  io_lineBuffer_o_data_55,
  output [7:0]  io_lineBuffer_o_data_56,
  output [7:0]  io_lineBuffer_o_data_57,
  output [7:0]  io_lineBuffer_o_data_58,
  output [7:0]  io_lineBuffer_o_data_59,
  output [7:0]  io_lineBuffer_o_data_60,
  output [7:0]  io_lineBuffer_o_data_61,
  output [7:0]  io_lineBuffer_o_data_62,
  output [7:0]  io_lineBuffer_o_data_63,
  output [7:0]  io_lineBuffer_o_data_64,
  output [7:0]  io_lineBuffer_o_data_65,
  output [7:0]  io_lineBuffer_o_data_66,
  output [7:0]  io_lineBuffer_o_data_67,
  output [7:0]  io_lineBuffer_o_data_68,
  output [7:0]  io_lineBuffer_o_data_69,
  output [7:0]  io_lineBuffer_o_data_70,
  output [7:0]  io_lineBuffer_o_data_71
);
  wire  buffer_0_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_0_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_0_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_0_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_0_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_0_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_1_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_1_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_1_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_1_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_1_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_1_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_2_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_2_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_2_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_2_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_2_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_2_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_3_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_3_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_3_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_3_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_3_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_3_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_4_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_4_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_4_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_4_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_4_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_4_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_5_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_5_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_5_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_5_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_5_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_5_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_6_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_6_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_6_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_6_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_6_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_6_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  wire  buffer_7_clock; // @[LineBuffer.scala 213:52]
  wire  buffer_7_reset; // @[LineBuffer.scala 213:52]
  wire [2:0] buffer_7_io_sel; // @[LineBuffer.scala 213:52]
  wire  buffer_7_io_s_mod; // @[LineBuffer.scala 213:52]
  wire [31:0] buffer_7_io_line_i_data; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_0; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_1; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_2; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_3; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_4; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_5; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_6; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_7; // @[LineBuffer.scala 213:52]
  wire [7:0] buffer_7_io_line_o_data_8; // @[LineBuffer.scala 213:52]
  line_buffer_unit_extend buffer_0 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_0_clock),
    .reset(buffer_0_reset),
    .io_sel(buffer_0_io_sel),
    .io_s_mod(buffer_0_io_s_mod),
    .io_line_i_data(buffer_0_io_line_i_data),
    .io_line_o_data_0(buffer_0_io_line_o_data_0),
    .io_line_o_data_1(buffer_0_io_line_o_data_1),
    .io_line_o_data_2(buffer_0_io_line_o_data_2),
    .io_line_o_data_3(buffer_0_io_line_o_data_3),
    .io_line_o_data_4(buffer_0_io_line_o_data_4),
    .io_line_o_data_5(buffer_0_io_line_o_data_5),
    .io_line_o_data_6(buffer_0_io_line_o_data_6),
    .io_line_o_data_7(buffer_0_io_line_o_data_7),
    .io_line_o_data_8(buffer_0_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_1 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_1_clock),
    .reset(buffer_1_reset),
    .io_sel(buffer_1_io_sel),
    .io_s_mod(buffer_1_io_s_mod),
    .io_line_i_data(buffer_1_io_line_i_data),
    .io_line_o_data_0(buffer_1_io_line_o_data_0),
    .io_line_o_data_1(buffer_1_io_line_o_data_1),
    .io_line_o_data_2(buffer_1_io_line_o_data_2),
    .io_line_o_data_3(buffer_1_io_line_o_data_3),
    .io_line_o_data_4(buffer_1_io_line_o_data_4),
    .io_line_o_data_5(buffer_1_io_line_o_data_5),
    .io_line_o_data_6(buffer_1_io_line_o_data_6),
    .io_line_o_data_7(buffer_1_io_line_o_data_7),
    .io_line_o_data_8(buffer_1_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_2 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_2_clock),
    .reset(buffer_2_reset),
    .io_sel(buffer_2_io_sel),
    .io_s_mod(buffer_2_io_s_mod),
    .io_line_i_data(buffer_2_io_line_i_data),
    .io_line_o_data_0(buffer_2_io_line_o_data_0),
    .io_line_o_data_1(buffer_2_io_line_o_data_1),
    .io_line_o_data_2(buffer_2_io_line_o_data_2),
    .io_line_o_data_3(buffer_2_io_line_o_data_3),
    .io_line_o_data_4(buffer_2_io_line_o_data_4),
    .io_line_o_data_5(buffer_2_io_line_o_data_5),
    .io_line_o_data_6(buffer_2_io_line_o_data_6),
    .io_line_o_data_7(buffer_2_io_line_o_data_7),
    .io_line_o_data_8(buffer_2_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_3 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_3_clock),
    .reset(buffer_3_reset),
    .io_sel(buffer_3_io_sel),
    .io_s_mod(buffer_3_io_s_mod),
    .io_line_i_data(buffer_3_io_line_i_data),
    .io_line_o_data_0(buffer_3_io_line_o_data_0),
    .io_line_o_data_1(buffer_3_io_line_o_data_1),
    .io_line_o_data_2(buffer_3_io_line_o_data_2),
    .io_line_o_data_3(buffer_3_io_line_o_data_3),
    .io_line_o_data_4(buffer_3_io_line_o_data_4),
    .io_line_o_data_5(buffer_3_io_line_o_data_5),
    .io_line_o_data_6(buffer_3_io_line_o_data_6),
    .io_line_o_data_7(buffer_3_io_line_o_data_7),
    .io_line_o_data_8(buffer_3_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_4 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_4_clock),
    .reset(buffer_4_reset),
    .io_sel(buffer_4_io_sel),
    .io_s_mod(buffer_4_io_s_mod),
    .io_line_i_data(buffer_4_io_line_i_data),
    .io_line_o_data_0(buffer_4_io_line_o_data_0),
    .io_line_o_data_1(buffer_4_io_line_o_data_1),
    .io_line_o_data_2(buffer_4_io_line_o_data_2),
    .io_line_o_data_3(buffer_4_io_line_o_data_3),
    .io_line_o_data_4(buffer_4_io_line_o_data_4),
    .io_line_o_data_5(buffer_4_io_line_o_data_5),
    .io_line_o_data_6(buffer_4_io_line_o_data_6),
    .io_line_o_data_7(buffer_4_io_line_o_data_7),
    .io_line_o_data_8(buffer_4_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_5 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_5_clock),
    .reset(buffer_5_reset),
    .io_sel(buffer_5_io_sel),
    .io_s_mod(buffer_5_io_s_mod),
    .io_line_i_data(buffer_5_io_line_i_data),
    .io_line_o_data_0(buffer_5_io_line_o_data_0),
    .io_line_o_data_1(buffer_5_io_line_o_data_1),
    .io_line_o_data_2(buffer_5_io_line_o_data_2),
    .io_line_o_data_3(buffer_5_io_line_o_data_3),
    .io_line_o_data_4(buffer_5_io_line_o_data_4),
    .io_line_o_data_5(buffer_5_io_line_o_data_5),
    .io_line_o_data_6(buffer_5_io_line_o_data_6),
    .io_line_o_data_7(buffer_5_io_line_o_data_7),
    .io_line_o_data_8(buffer_5_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_6 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_6_clock),
    .reset(buffer_6_reset),
    .io_sel(buffer_6_io_sel),
    .io_s_mod(buffer_6_io_s_mod),
    .io_line_i_data(buffer_6_io_line_i_data),
    .io_line_o_data_0(buffer_6_io_line_o_data_0),
    .io_line_o_data_1(buffer_6_io_line_o_data_1),
    .io_line_o_data_2(buffer_6_io_line_o_data_2),
    .io_line_o_data_3(buffer_6_io_line_o_data_3),
    .io_line_o_data_4(buffer_6_io_line_o_data_4),
    .io_line_o_data_5(buffer_6_io_line_o_data_5),
    .io_line_o_data_6(buffer_6_io_line_o_data_6),
    .io_line_o_data_7(buffer_6_io_line_o_data_7),
    .io_line_o_data_8(buffer_6_io_line_o_data_8)
  );
  line_buffer_unit_extend buffer_7 ( // @[LineBuffer.scala 213:52]
    .clock(buffer_7_clock),
    .reset(buffer_7_reset),
    .io_sel(buffer_7_io_sel),
    .io_s_mod(buffer_7_io_s_mod),
    .io_line_i_data(buffer_7_io_line_i_data),
    .io_line_o_data_0(buffer_7_io_line_o_data_0),
    .io_line_o_data_1(buffer_7_io_line_o_data_1),
    .io_line_o_data_2(buffer_7_io_line_o_data_2),
    .io_line_o_data_3(buffer_7_io_line_o_data_3),
    .io_line_o_data_4(buffer_7_io_line_o_data_4),
    .io_line_o_data_5(buffer_7_io_line_o_data_5),
    .io_line_o_data_6(buffer_7_io_line_o_data_6),
    .io_line_o_data_7(buffer_7_io_line_o_data_7),
    .io_line_o_data_8(buffer_7_io_line_o_data_8)
  );
  assign io_lineBuffer_o_data_0 = buffer_0_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_1 = buffer_0_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_2 = buffer_0_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_3 = buffer_0_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_4 = buffer_0_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_5 = buffer_0_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_6 = buffer_0_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_7 = buffer_0_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_8 = buffer_0_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_9 = buffer_1_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_10 = buffer_1_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_11 = buffer_1_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_12 = buffer_1_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_13 = buffer_1_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_14 = buffer_1_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_15 = buffer_1_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_16 = buffer_1_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_17 = buffer_1_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_18 = buffer_2_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_19 = buffer_2_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_20 = buffer_2_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_21 = buffer_2_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_22 = buffer_2_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_23 = buffer_2_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_24 = buffer_2_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_25 = buffer_2_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_26 = buffer_2_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_27 = buffer_3_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_28 = buffer_3_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_29 = buffer_3_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_30 = buffer_3_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_31 = buffer_3_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_32 = buffer_3_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_33 = buffer_3_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_34 = buffer_3_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_35 = buffer_3_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_36 = buffer_4_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_37 = buffer_4_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_38 = buffer_4_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_39 = buffer_4_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_40 = buffer_4_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_41 = buffer_4_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_42 = buffer_4_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_43 = buffer_4_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_44 = buffer_4_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_45 = buffer_5_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_46 = buffer_5_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_47 = buffer_5_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_48 = buffer_5_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_49 = buffer_5_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_50 = buffer_5_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_51 = buffer_5_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_52 = buffer_5_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_53 = buffer_5_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_54 = buffer_6_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_55 = buffer_6_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_56 = buffer_6_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_57 = buffer_6_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_58 = buffer_6_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_59 = buffer_6_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_60 = buffer_6_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_61 = buffer_6_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_62 = buffer_6_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_63 = buffer_7_io_line_o_data_0; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_64 = buffer_7_io_line_o_data_1; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_65 = buffer_7_io_line_o_data_2; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_66 = buffer_7_io_line_o_data_3; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_67 = buffer_7_io_line_o_data_4; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_68 = buffer_7_io_line_o_data_5; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_69 = buffer_7_io_line_o_data_6; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_70 = buffer_7_io_line_o_data_7; // @[LineBuffer.scala 221:45]
  assign io_lineBuffer_o_data_71 = buffer_7_io_line_o_data_8; // @[LineBuffer.scala 221:45]
  assign buffer_0_clock = clock;
  assign buffer_0_reset = reset;
  assign buffer_0_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_0_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_0_io_line_i_data = io_lineBuffer_i_data_0; // @[LineBuffer.scala 219:34]
  assign buffer_1_clock = clock;
  assign buffer_1_reset = reset;
  assign buffer_1_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_1_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_1_io_line_i_data = io_lineBuffer_i_data_1; // @[LineBuffer.scala 219:34]
  assign buffer_2_clock = clock;
  assign buffer_2_reset = reset;
  assign buffer_2_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_2_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_2_io_line_i_data = io_lineBuffer_i_data_2; // @[LineBuffer.scala 219:34]
  assign buffer_3_clock = clock;
  assign buffer_3_reset = reset;
  assign buffer_3_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_3_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_3_io_line_i_data = io_lineBuffer_i_data_3; // @[LineBuffer.scala 219:34]
  assign buffer_4_clock = clock;
  assign buffer_4_reset = reset;
  assign buffer_4_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_4_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_4_io_line_i_data = io_lineBuffer_i_data_4; // @[LineBuffer.scala 219:34]
  assign buffer_5_clock = clock;
  assign buffer_5_reset = reset;
  assign buffer_5_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_5_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_5_io_line_i_data = io_lineBuffer_i_data_5; // @[LineBuffer.scala 219:34]
  assign buffer_6_clock = clock;
  assign buffer_6_reset = reset;
  assign buffer_6_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_6_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_6_io_line_i_data = io_lineBuffer_i_data_6; // @[LineBuffer.scala 219:34]
  assign buffer_7_clock = clock;
  assign buffer_7_reset = reset;
  assign buffer_7_io_sel = io_sel; // @[LineBuffer.scala 215:26]
  assign buffer_7_io_s_mod = io_s_mod; // @[LineBuffer.scala 217:28]
  assign buffer_7_io_line_i_data = io_lineBuffer_i_data_7; // @[LineBuffer.scala 219:34]
endmodule
module mult_int8_2(
  input         clock,
  input  [7:0]  io_a,
  input  [7:0]  io_b,
  input  [7:0]  io_c,
  output [15:0] io_ac,
  output [15:0] io_bc
);
  wire  cal_mult_clk; // @[utils.scala 624:26]
  wire [7:0] cal_mult_a; // @[utils.scala 624:26]
  wire [7:0] cal_mult_b; // @[utils.scala 624:26]
  wire [7:0] cal_mult_c; // @[utils.scala 624:26]
  wire [15:0] cal_mult_ac; // @[utils.scala 624:26]
  wire [15:0] cal_mult_bc; // @[utils.scala 624:26]
  wire [15:0] bc_temp = cal_mult_bc; // @[utils.scala 622:23 629:13]
  wire [15:0] _GEN_0 = {{15'd0}, bc_temp[15]}; // @[utils.scala 631:32]
  wire [15:0] ac_temp = cal_mult_ac; // @[utils.scala 621:23 628:13]
  wire [15:0] _ac_comp_T_4 = $signed(ac_temp) + 16'sh1; // @[utils.scala 631:55]
  cal_mult_int8_x2_dsp cal_mult ( // @[utils.scala 624:26]
    .clk(cal_mult_clk),
    .a(cal_mult_a),
    .b(cal_mult_b),
    .c(cal_mult_c),
    .ac(cal_mult_ac),
    .bc(cal_mult_bc)
  );
  assign io_ac = _GEN_0 == 16'h1 ? $signed(_ac_comp_T_4) : $signed(ac_temp); // @[utils.scala 631:19]
  assign io_bc = cal_mult_bc; // @[utils.scala 622:23 629:13]
  assign cal_mult_clk = clock; // @[utils.scala 630:21]
  assign cal_mult_a = io_a; // @[utils.scala 625:19]
  assign cal_mult_b = io_b; // @[utils.scala 626:19]
  assign cal_mult_c = io_c; // @[utils.scala 627:19]
endmodule
module addtree_int16_3_3(
  input         clock,
  input  [15:0] io_din_0,
  input  [15:0] io_din_1,
  input  [15:0] io_din_2,
  input  [15:0] io_din_3,
  input  [15:0] io_din_4,
  input  [15:0] io_din_5,
  input  [15:0] io_din_6,
  input  [15:0] io_din_7,
  input  [15:0] io_din_8,
  output [17:0] io_dout
);
  wire  addtree_clk; // @[utils.scala 662:25]
  wire [15:0] addtree_a1; // @[utils.scala 662:25]
  wire [15:0] addtree_a2; // @[utils.scala 662:25]
  wire [15:0] addtree_a3; // @[utils.scala 662:25]
  wire [15:0] addtree_a4; // @[utils.scala 662:25]
  wire [15:0] addtree_a5; // @[utils.scala 662:25]
  wire [15:0] addtree_a6; // @[utils.scala 662:25]
  wire [15:0] addtree_a7; // @[utils.scala 662:25]
  wire [15:0] addtree_a8; // @[utils.scala 662:25]
  wire [15:0] addtree_a9; // @[utils.scala 662:25]
  wire [17:0] addtree_dout; // @[utils.scala 662:25]
  cal_addtree_int16_x9 addtree ( // @[utils.scala 662:25]
    .clk(addtree_clk),
    .a1(addtree_a1),
    .a2(addtree_a2),
    .a3(addtree_a3),
    .a4(addtree_a4),
    .a5(addtree_a5),
    .a6(addtree_a6),
    .a7(addtree_a7),
    .a8(addtree_a8),
    .a9(addtree_a9),
    .dout(addtree_dout)
  );
  assign io_dout = addtree_dout; // @[utils.scala 673:13]
  assign addtree_clk = clock; // @[utils.scala 663:20]
  assign addtree_a1 = io_din_0; // @[utils.scala 664:19]
  assign addtree_a2 = io_din_1; // @[utils.scala 665:19]
  assign addtree_a3 = io_din_2; // @[utils.scala 666:19]
  assign addtree_a4 = io_din_3; // @[utils.scala 667:19]
  assign addtree_a5 = io_din_4; // @[utils.scala 668:19]
  assign addtree_a6 = io_din_5; // @[utils.scala 669:19]
  assign addtree_a7 = io_din_6; // @[utils.scala 670:19]
  assign addtree_a8 = io_din_7; // @[utils.scala 671:19]
  assign addtree_a9 = io_din_8; // @[utils.scala 672:19]
endmodule
module conv_win_3_3(
  input         clock,
  input  [7:0]  io_ifm_win_33_0,
  input  [7:0]  io_ifm_win_33_1,
  input  [7:0]  io_ifm_win_33_2,
  input  [7:0]  io_ifm_win_33_3,
  input  [7:0]  io_ifm_win_33_4,
  input  [7:0]  io_ifm_win_33_5,
  input  [7:0]  io_ifm_win_33_6,
  input  [7:0]  io_ifm_win_33_7,
  input  [7:0]  io_ifm_win_33_8,
  input  [7:0]  io_weight_win_33_ch1_0,
  input  [7:0]  io_weight_win_33_ch1_1,
  input  [7:0]  io_weight_win_33_ch1_2,
  input  [7:0]  io_weight_win_33_ch1_3,
  input  [7:0]  io_weight_win_33_ch1_4,
  input  [7:0]  io_weight_win_33_ch1_5,
  input  [7:0]  io_weight_win_33_ch1_6,
  input  [7:0]  io_weight_win_33_ch1_7,
  input  [7:0]  io_weight_win_33_ch1_8,
  input  [7:0]  io_weight_win_33_ch2_0,
  input  [7:0]  io_weight_win_33_ch2_1,
  input  [7:0]  io_weight_win_33_ch2_2,
  input  [7:0]  io_weight_win_33_ch2_3,
  input  [7:0]  io_weight_win_33_ch2_4,
  input  [7:0]  io_weight_win_33_ch2_5,
  input  [7:0]  io_weight_win_33_ch2_6,
  input  [7:0]  io_weight_win_33_ch2_7,
  input  [7:0]  io_weight_win_33_ch2_8,
  output [17:0] io_o_conv_ch1,
  output [17:0] io_o_conv_ch2
);
  wire  mult_0_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_0_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_0_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_0_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_0_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_0_io_bc; // @[Conv.scala 83:34]
  wire  mult_1_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_1_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_1_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_1_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_1_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_1_io_bc; // @[Conv.scala 83:34]
  wire  mult_2_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_2_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_2_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_2_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_2_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_2_io_bc; // @[Conv.scala 83:34]
  wire  mult_3_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_3_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_3_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_3_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_3_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_3_io_bc; // @[Conv.scala 83:34]
  wire  mult_4_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_4_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_4_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_4_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_4_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_4_io_bc; // @[Conv.scala 83:34]
  wire  mult_5_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_5_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_5_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_5_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_5_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_5_io_bc; // @[Conv.scala 83:34]
  wire  mult_6_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_6_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_6_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_6_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_6_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_6_io_bc; // @[Conv.scala 83:34]
  wire  mult_7_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_7_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_7_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_7_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_7_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_7_io_bc; // @[Conv.scala 83:34]
  wire  mult_8_clock; // @[Conv.scala 83:34]
  wire [7:0] mult_8_io_a; // @[Conv.scala 83:34]
  wire [7:0] mult_8_io_b; // @[Conv.scala 83:34]
  wire [7:0] mult_8_io_c; // @[Conv.scala 83:34]
  wire [15:0] mult_8_io_ac; // @[Conv.scala 83:34]
  wire [15:0] mult_8_io_bc; // @[Conv.scala 83:34]
  wire  addtree_0_clock; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_0; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_1; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_2; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_3; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_4; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_5; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_6; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_7; // @[Conv.scala 92:37]
  wire [15:0] addtree_0_io_din_8; // @[Conv.scala 92:37]
  wire [17:0] addtree_0_io_dout; // @[Conv.scala 92:37]
  wire  addtree_1_clock; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_0; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_1; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_2; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_3; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_4; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_5; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_6; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_7; // @[Conv.scala 92:37]
  wire [15:0] addtree_1_io_din_8; // @[Conv.scala 92:37]
  wire [17:0] addtree_1_io_dout; // @[Conv.scala 92:37]
  mult_int8_2 mult_0 ( // @[Conv.scala 83:34]
    .clock(mult_0_clock),
    .io_a(mult_0_io_a),
    .io_b(mult_0_io_b),
    .io_c(mult_0_io_c),
    .io_ac(mult_0_io_ac),
    .io_bc(mult_0_io_bc)
  );
  mult_int8_2 mult_1 ( // @[Conv.scala 83:34]
    .clock(mult_1_clock),
    .io_a(mult_1_io_a),
    .io_b(mult_1_io_b),
    .io_c(mult_1_io_c),
    .io_ac(mult_1_io_ac),
    .io_bc(mult_1_io_bc)
  );
  mult_int8_2 mult_2 ( // @[Conv.scala 83:34]
    .clock(mult_2_clock),
    .io_a(mult_2_io_a),
    .io_b(mult_2_io_b),
    .io_c(mult_2_io_c),
    .io_ac(mult_2_io_ac),
    .io_bc(mult_2_io_bc)
  );
  mult_int8_2 mult_3 ( // @[Conv.scala 83:34]
    .clock(mult_3_clock),
    .io_a(mult_3_io_a),
    .io_b(mult_3_io_b),
    .io_c(mult_3_io_c),
    .io_ac(mult_3_io_ac),
    .io_bc(mult_3_io_bc)
  );
  mult_int8_2 mult_4 ( // @[Conv.scala 83:34]
    .clock(mult_4_clock),
    .io_a(mult_4_io_a),
    .io_b(mult_4_io_b),
    .io_c(mult_4_io_c),
    .io_ac(mult_4_io_ac),
    .io_bc(mult_4_io_bc)
  );
  mult_int8_2 mult_5 ( // @[Conv.scala 83:34]
    .clock(mult_5_clock),
    .io_a(mult_5_io_a),
    .io_b(mult_5_io_b),
    .io_c(mult_5_io_c),
    .io_ac(mult_5_io_ac),
    .io_bc(mult_5_io_bc)
  );
  mult_int8_2 mult_6 ( // @[Conv.scala 83:34]
    .clock(mult_6_clock),
    .io_a(mult_6_io_a),
    .io_b(mult_6_io_b),
    .io_c(mult_6_io_c),
    .io_ac(mult_6_io_ac),
    .io_bc(mult_6_io_bc)
  );
  mult_int8_2 mult_7 ( // @[Conv.scala 83:34]
    .clock(mult_7_clock),
    .io_a(mult_7_io_a),
    .io_b(mult_7_io_b),
    .io_c(mult_7_io_c),
    .io_ac(mult_7_io_ac),
    .io_bc(mult_7_io_bc)
  );
  mult_int8_2 mult_8 ( // @[Conv.scala 83:34]
    .clock(mult_8_clock),
    .io_a(mult_8_io_a),
    .io_b(mult_8_io_b),
    .io_c(mult_8_io_c),
    .io_ac(mult_8_io_ac),
    .io_bc(mult_8_io_bc)
  );
  addtree_int16_3_3 addtree_0 ( // @[Conv.scala 92:37]
    .clock(addtree_0_clock),
    .io_din_0(addtree_0_io_din_0),
    .io_din_1(addtree_0_io_din_1),
    .io_din_2(addtree_0_io_din_2),
    .io_din_3(addtree_0_io_din_3),
    .io_din_4(addtree_0_io_din_4),
    .io_din_5(addtree_0_io_din_5),
    .io_din_6(addtree_0_io_din_6),
    .io_din_7(addtree_0_io_din_7),
    .io_din_8(addtree_0_io_din_8),
    .io_dout(addtree_0_io_dout)
  );
  addtree_int16_3_3 addtree_1 ( // @[Conv.scala 92:37]
    .clock(addtree_1_clock),
    .io_din_0(addtree_1_io_din_0),
    .io_din_1(addtree_1_io_din_1),
    .io_din_2(addtree_1_io_din_2),
    .io_din_3(addtree_1_io_din_3),
    .io_din_4(addtree_1_io_din_4),
    .io_din_5(addtree_1_io_din_5),
    .io_din_6(addtree_1_io_din_6),
    .io_din_7(addtree_1_io_din_7),
    .io_din_8(addtree_1_io_din_8),
    .io_dout(addtree_1_io_dout)
  );
  assign io_o_conv_ch1 = addtree_0_io_dout; // @[Conv.scala 97:41]
  assign io_o_conv_ch2 = addtree_1_io_dout; // @[Conv.scala 98:41]
  assign mult_0_clock = clock;
  assign mult_0_io_a = io_weight_win_33_ch1_0; // @[Conv.scala 86:49]
  assign mult_0_io_b = io_weight_win_33_ch2_0; // @[Conv.scala 87:49]
  assign mult_0_io_c = io_ifm_win_33_0; // @[Conv.scala 85:42]
  assign mult_1_clock = clock;
  assign mult_1_io_a = io_weight_win_33_ch1_1; // @[Conv.scala 86:49]
  assign mult_1_io_b = io_weight_win_33_ch2_1; // @[Conv.scala 87:49]
  assign mult_1_io_c = io_ifm_win_33_1; // @[Conv.scala 85:42]
  assign mult_2_clock = clock;
  assign mult_2_io_a = io_weight_win_33_ch1_2; // @[Conv.scala 86:49]
  assign mult_2_io_b = io_weight_win_33_ch2_2; // @[Conv.scala 87:49]
  assign mult_2_io_c = io_ifm_win_33_2; // @[Conv.scala 85:42]
  assign mult_3_clock = clock;
  assign mult_3_io_a = io_weight_win_33_ch1_3; // @[Conv.scala 86:49]
  assign mult_3_io_b = io_weight_win_33_ch2_3; // @[Conv.scala 87:49]
  assign mult_3_io_c = io_ifm_win_33_3; // @[Conv.scala 85:42]
  assign mult_4_clock = clock;
  assign mult_4_io_a = io_weight_win_33_ch1_4; // @[Conv.scala 86:49]
  assign mult_4_io_b = io_weight_win_33_ch2_4; // @[Conv.scala 87:49]
  assign mult_4_io_c = io_ifm_win_33_4; // @[Conv.scala 85:42]
  assign mult_5_clock = clock;
  assign mult_5_io_a = io_weight_win_33_ch1_5; // @[Conv.scala 86:49]
  assign mult_5_io_b = io_weight_win_33_ch2_5; // @[Conv.scala 87:49]
  assign mult_5_io_c = io_ifm_win_33_5; // @[Conv.scala 85:42]
  assign mult_6_clock = clock;
  assign mult_6_io_a = io_weight_win_33_ch1_6; // @[Conv.scala 86:49]
  assign mult_6_io_b = io_weight_win_33_ch2_6; // @[Conv.scala 87:49]
  assign mult_6_io_c = io_ifm_win_33_6; // @[Conv.scala 85:42]
  assign mult_7_clock = clock;
  assign mult_7_io_a = io_weight_win_33_ch1_7; // @[Conv.scala 86:49]
  assign mult_7_io_b = io_weight_win_33_ch2_7; // @[Conv.scala 87:49]
  assign mult_7_io_c = io_ifm_win_33_7; // @[Conv.scala 85:42]
  assign mult_8_clock = clock;
  assign mult_8_io_a = io_weight_win_33_ch1_8; // @[Conv.scala 86:49]
  assign mult_8_io_b = io_weight_win_33_ch2_8; // @[Conv.scala 87:49]
  assign mult_8_io_c = io_ifm_win_33_8; // @[Conv.scala 85:42]
  assign addtree_0_clock = clock;
  assign addtree_0_io_din_0 = mult_0_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_1 = mult_1_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_2 = mult_2_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_3 = mult_3_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_4 = mult_4_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_5 = mult_5_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_6 = mult_6_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_7 = mult_7_io_ac; // @[Conv.scala 94:40]
  assign addtree_0_io_din_8 = mult_8_io_ac; // @[Conv.scala 94:40]
  assign addtree_1_clock = clock;
  assign addtree_1_io_din_0 = mult_0_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_1 = mult_1_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_2 = mult_2_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_3 = mult_3_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_4 = mult_4_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_5 = mult_5_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_6 = mult_6_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_7 = mult_7_io_bc; // @[Conv.scala 95:40]
  assign addtree_1_io_din_8 = mult_8_io_bc; // @[Conv.scala 95:40]
endmodule
module addtree_int18_3_3(
  input         clock,
  input  [17:0] io_din_0,
  input  [17:0] io_din_1,
  input  [17:0] io_din_2,
  input  [17:0] io_din_3,
  input  [17:0] io_din_4,
  input  [17:0] io_din_5,
  input  [17:0] io_din_6,
  input  [17:0] io_din_7,
  input  [17:0] io_bias,
  output [17:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] temp_0; // @[utils.scala 707:19]
  reg [17:0] temp_1; // @[utils.scala 707:19]
  reg [17:0] temp_2; // @[utils.scala 707:19]
  reg [17:0] temp_3; // @[utils.scala 707:19]
  wire [17:0] _temp_0_T_2 = $signed(io_din_0) + $signed(io_din_1); // @[utils.scala 708:22]
  wire [17:0] _temp_1_T_2 = $signed(io_din_3) + $signed(io_din_4); // @[utils.scala 709:22]
  wire [17:0] _temp_2_T_2 = $signed(io_din_6) + $signed(io_din_7); // @[utils.scala 710:22]
  wire [17:0] _temp_3_T_2 = $signed(temp_0) + $signed(temp_1); // @[utils.scala 711:24]
  assign io_dout = temp_3; // @[utils.scala 712:24]
  always @(posedge clock) begin
    temp_0 <= $signed(_temp_0_T_2) + $signed(io_din_2); // @[utils.scala 708:30]
    temp_1 <= $signed(_temp_1_T_2) + $signed(io_din_5); // @[utils.scala 709:30]
    temp_2 <= $signed(_temp_2_T_2) + $signed(io_bias); // @[utils.scala 710:30]
    temp_3 <= $signed(_temp_3_T_2) + $signed(temp_2); // @[utils.scala 711:34]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  temp_1 = _RAND_1[17:0];
  _RAND_2 = {1{`RANDOM}};
  temp_2 = _RAND_2[17:0];
  _RAND_3 = {1{`RANDOM}};
  temp_3 = _RAND_3[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module conv_unit(
  input         clock,
  input  [7:0]  io_ifm_win_33_0,
  input  [7:0]  io_ifm_win_33_1,
  input  [7:0]  io_ifm_win_33_2,
  input  [7:0]  io_ifm_win_33_3,
  input  [7:0]  io_ifm_win_33_4,
  input  [7:0]  io_ifm_win_33_5,
  input  [7:0]  io_ifm_win_33_6,
  input  [7:0]  io_ifm_win_33_7,
  input  [7:0]  io_ifm_win_33_8,
  input  [7:0]  io_ifm_win_33_9,
  input  [7:0]  io_ifm_win_33_10,
  input  [7:0]  io_ifm_win_33_11,
  input  [7:0]  io_ifm_win_33_12,
  input  [7:0]  io_ifm_win_33_13,
  input  [7:0]  io_ifm_win_33_14,
  input  [7:0]  io_ifm_win_33_15,
  input  [7:0]  io_ifm_win_33_16,
  input  [7:0]  io_ifm_win_33_17,
  input  [7:0]  io_ifm_win_33_18,
  input  [7:0]  io_ifm_win_33_19,
  input  [7:0]  io_ifm_win_33_20,
  input  [7:0]  io_ifm_win_33_21,
  input  [7:0]  io_ifm_win_33_22,
  input  [7:0]  io_ifm_win_33_23,
  input  [7:0]  io_ifm_win_33_24,
  input  [7:0]  io_ifm_win_33_25,
  input  [7:0]  io_ifm_win_33_26,
  input  [7:0]  io_ifm_win_33_27,
  input  [7:0]  io_ifm_win_33_28,
  input  [7:0]  io_ifm_win_33_29,
  input  [7:0]  io_ifm_win_33_30,
  input  [7:0]  io_ifm_win_33_31,
  input  [7:0]  io_ifm_win_33_32,
  input  [7:0]  io_ifm_win_33_33,
  input  [7:0]  io_ifm_win_33_34,
  input  [7:0]  io_ifm_win_33_35,
  input  [7:0]  io_ifm_win_33_36,
  input  [7:0]  io_ifm_win_33_37,
  input  [7:0]  io_ifm_win_33_38,
  input  [7:0]  io_ifm_win_33_39,
  input  [7:0]  io_ifm_win_33_40,
  input  [7:0]  io_ifm_win_33_41,
  input  [7:0]  io_ifm_win_33_42,
  input  [7:0]  io_ifm_win_33_43,
  input  [7:0]  io_ifm_win_33_44,
  input  [7:0]  io_ifm_win_33_45,
  input  [7:0]  io_ifm_win_33_46,
  input  [7:0]  io_ifm_win_33_47,
  input  [7:0]  io_ifm_win_33_48,
  input  [7:0]  io_ifm_win_33_49,
  input  [7:0]  io_ifm_win_33_50,
  input  [7:0]  io_ifm_win_33_51,
  input  [7:0]  io_ifm_win_33_52,
  input  [7:0]  io_ifm_win_33_53,
  input  [7:0]  io_ifm_win_33_54,
  input  [7:0]  io_ifm_win_33_55,
  input  [7:0]  io_ifm_win_33_56,
  input  [7:0]  io_ifm_win_33_57,
  input  [7:0]  io_ifm_win_33_58,
  input  [7:0]  io_ifm_win_33_59,
  input  [7:0]  io_ifm_win_33_60,
  input  [7:0]  io_ifm_win_33_61,
  input  [7:0]  io_ifm_win_33_62,
  input  [7:0]  io_ifm_win_33_63,
  input  [7:0]  io_ifm_win_33_64,
  input  [7:0]  io_ifm_win_33_65,
  input  [7:0]  io_ifm_win_33_66,
  input  [7:0]  io_ifm_win_33_67,
  input  [7:0]  io_ifm_win_33_68,
  input  [7:0]  io_ifm_win_33_69,
  input  [7:0]  io_ifm_win_33_70,
  input  [7:0]  io_ifm_win_33_71,
  input  [7:0]  io_weight_win_33_ch1_0,
  input  [7:0]  io_weight_win_33_ch1_1,
  input  [7:0]  io_weight_win_33_ch1_2,
  input  [7:0]  io_weight_win_33_ch1_3,
  input  [7:0]  io_weight_win_33_ch1_4,
  input  [7:0]  io_weight_win_33_ch1_5,
  input  [7:0]  io_weight_win_33_ch1_6,
  input  [7:0]  io_weight_win_33_ch1_7,
  input  [7:0]  io_weight_win_33_ch1_8,
  input  [7:0]  io_weight_win_33_ch1_9,
  input  [7:0]  io_weight_win_33_ch1_10,
  input  [7:0]  io_weight_win_33_ch1_11,
  input  [7:0]  io_weight_win_33_ch1_12,
  input  [7:0]  io_weight_win_33_ch1_13,
  input  [7:0]  io_weight_win_33_ch1_14,
  input  [7:0]  io_weight_win_33_ch1_15,
  input  [7:0]  io_weight_win_33_ch1_16,
  input  [7:0]  io_weight_win_33_ch1_17,
  input  [7:0]  io_weight_win_33_ch1_18,
  input  [7:0]  io_weight_win_33_ch1_19,
  input  [7:0]  io_weight_win_33_ch1_20,
  input  [7:0]  io_weight_win_33_ch1_21,
  input  [7:0]  io_weight_win_33_ch1_22,
  input  [7:0]  io_weight_win_33_ch1_23,
  input  [7:0]  io_weight_win_33_ch1_24,
  input  [7:0]  io_weight_win_33_ch1_25,
  input  [7:0]  io_weight_win_33_ch1_26,
  input  [7:0]  io_weight_win_33_ch1_27,
  input  [7:0]  io_weight_win_33_ch1_28,
  input  [7:0]  io_weight_win_33_ch1_29,
  input  [7:0]  io_weight_win_33_ch1_30,
  input  [7:0]  io_weight_win_33_ch1_31,
  input  [7:0]  io_weight_win_33_ch1_32,
  input  [7:0]  io_weight_win_33_ch1_33,
  input  [7:0]  io_weight_win_33_ch1_34,
  input  [7:0]  io_weight_win_33_ch1_35,
  input  [7:0]  io_weight_win_33_ch1_36,
  input  [7:0]  io_weight_win_33_ch1_37,
  input  [7:0]  io_weight_win_33_ch1_38,
  input  [7:0]  io_weight_win_33_ch1_39,
  input  [7:0]  io_weight_win_33_ch1_40,
  input  [7:0]  io_weight_win_33_ch1_41,
  input  [7:0]  io_weight_win_33_ch1_42,
  input  [7:0]  io_weight_win_33_ch1_43,
  input  [7:0]  io_weight_win_33_ch1_44,
  input  [7:0]  io_weight_win_33_ch1_45,
  input  [7:0]  io_weight_win_33_ch1_46,
  input  [7:0]  io_weight_win_33_ch1_47,
  input  [7:0]  io_weight_win_33_ch1_48,
  input  [7:0]  io_weight_win_33_ch1_49,
  input  [7:0]  io_weight_win_33_ch1_50,
  input  [7:0]  io_weight_win_33_ch1_51,
  input  [7:0]  io_weight_win_33_ch1_52,
  input  [7:0]  io_weight_win_33_ch1_53,
  input  [7:0]  io_weight_win_33_ch1_54,
  input  [7:0]  io_weight_win_33_ch1_55,
  input  [7:0]  io_weight_win_33_ch1_56,
  input  [7:0]  io_weight_win_33_ch1_57,
  input  [7:0]  io_weight_win_33_ch1_58,
  input  [7:0]  io_weight_win_33_ch1_59,
  input  [7:0]  io_weight_win_33_ch1_60,
  input  [7:0]  io_weight_win_33_ch1_61,
  input  [7:0]  io_weight_win_33_ch1_62,
  input  [7:0]  io_weight_win_33_ch1_63,
  input  [7:0]  io_weight_win_33_ch1_64,
  input  [7:0]  io_weight_win_33_ch1_65,
  input  [7:0]  io_weight_win_33_ch1_66,
  input  [7:0]  io_weight_win_33_ch1_67,
  input  [7:0]  io_weight_win_33_ch1_68,
  input  [7:0]  io_weight_win_33_ch1_69,
  input  [7:0]  io_weight_win_33_ch1_70,
  input  [7:0]  io_weight_win_33_ch1_71,
  input  [7:0]  io_weight_win_33_ch2_0,
  input  [7:0]  io_weight_win_33_ch2_1,
  input  [7:0]  io_weight_win_33_ch2_2,
  input  [7:0]  io_weight_win_33_ch2_3,
  input  [7:0]  io_weight_win_33_ch2_4,
  input  [7:0]  io_weight_win_33_ch2_5,
  input  [7:0]  io_weight_win_33_ch2_6,
  input  [7:0]  io_weight_win_33_ch2_7,
  input  [7:0]  io_weight_win_33_ch2_8,
  input  [7:0]  io_weight_win_33_ch2_9,
  input  [7:0]  io_weight_win_33_ch2_10,
  input  [7:0]  io_weight_win_33_ch2_11,
  input  [7:0]  io_weight_win_33_ch2_12,
  input  [7:0]  io_weight_win_33_ch2_13,
  input  [7:0]  io_weight_win_33_ch2_14,
  input  [7:0]  io_weight_win_33_ch2_15,
  input  [7:0]  io_weight_win_33_ch2_16,
  input  [7:0]  io_weight_win_33_ch2_17,
  input  [7:0]  io_weight_win_33_ch2_18,
  input  [7:0]  io_weight_win_33_ch2_19,
  input  [7:0]  io_weight_win_33_ch2_20,
  input  [7:0]  io_weight_win_33_ch2_21,
  input  [7:0]  io_weight_win_33_ch2_22,
  input  [7:0]  io_weight_win_33_ch2_23,
  input  [7:0]  io_weight_win_33_ch2_24,
  input  [7:0]  io_weight_win_33_ch2_25,
  input  [7:0]  io_weight_win_33_ch2_26,
  input  [7:0]  io_weight_win_33_ch2_27,
  input  [7:0]  io_weight_win_33_ch2_28,
  input  [7:0]  io_weight_win_33_ch2_29,
  input  [7:0]  io_weight_win_33_ch2_30,
  input  [7:0]  io_weight_win_33_ch2_31,
  input  [7:0]  io_weight_win_33_ch2_32,
  input  [7:0]  io_weight_win_33_ch2_33,
  input  [7:0]  io_weight_win_33_ch2_34,
  input  [7:0]  io_weight_win_33_ch2_35,
  input  [7:0]  io_weight_win_33_ch2_36,
  input  [7:0]  io_weight_win_33_ch2_37,
  input  [7:0]  io_weight_win_33_ch2_38,
  input  [7:0]  io_weight_win_33_ch2_39,
  input  [7:0]  io_weight_win_33_ch2_40,
  input  [7:0]  io_weight_win_33_ch2_41,
  input  [7:0]  io_weight_win_33_ch2_42,
  input  [7:0]  io_weight_win_33_ch2_43,
  input  [7:0]  io_weight_win_33_ch2_44,
  input  [7:0]  io_weight_win_33_ch2_45,
  input  [7:0]  io_weight_win_33_ch2_46,
  input  [7:0]  io_weight_win_33_ch2_47,
  input  [7:0]  io_weight_win_33_ch2_48,
  input  [7:0]  io_weight_win_33_ch2_49,
  input  [7:0]  io_weight_win_33_ch2_50,
  input  [7:0]  io_weight_win_33_ch2_51,
  input  [7:0]  io_weight_win_33_ch2_52,
  input  [7:0]  io_weight_win_33_ch2_53,
  input  [7:0]  io_weight_win_33_ch2_54,
  input  [7:0]  io_weight_win_33_ch2_55,
  input  [7:0]  io_weight_win_33_ch2_56,
  input  [7:0]  io_weight_win_33_ch2_57,
  input  [7:0]  io_weight_win_33_ch2_58,
  input  [7:0]  io_weight_win_33_ch2_59,
  input  [7:0]  io_weight_win_33_ch2_60,
  input  [7:0]  io_weight_win_33_ch2_61,
  input  [7:0]  io_weight_win_33_ch2_62,
  input  [7:0]  io_weight_win_33_ch2_63,
  input  [7:0]  io_weight_win_33_ch2_64,
  input  [7:0]  io_weight_win_33_ch2_65,
  input  [7:0]  io_weight_win_33_ch2_66,
  input  [7:0]  io_weight_win_33_ch2_67,
  input  [7:0]  io_weight_win_33_ch2_68,
  input  [7:0]  io_weight_win_33_ch2_69,
  input  [7:0]  io_weight_win_33_ch2_70,
  input  [7:0]  io_weight_win_33_ch2_71,
  input  [17:0] io_bias1,
  input  [17:0] io_bias2,
  input         io_bias_valid,
  output [17:0] io_o_conv_ch1,
  output [17:0] io_o_conv_ch2
);
  wire  conv_33_0_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_0_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_0_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_0_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_1_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_1_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_1_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_1_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_2_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_2_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_2_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_2_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_3_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_3_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_3_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_3_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_4_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_4_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_4_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_4_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_5_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_5_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_5_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_5_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_6_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_6_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_6_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_6_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  conv_33_7_clock; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_ifm_win_33_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch1_8; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_0; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_1; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_2; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_3; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_4; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_5; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_6; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_7; // @[Conv.scala 47:40]
  wire [7:0] conv_33_7_io_weight_win_33_ch2_8; // @[Conv.scala 47:40]
  wire [17:0] conv_33_7_io_o_conv_ch1; // @[Conv.scala 47:40]
  wire [17:0] conv_33_7_io_o_conv_ch2; // @[Conv.scala 47:40]
  wire  addtree_0_clock; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_0; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_1; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_2; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_3; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_4; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_5; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_6; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_din_7; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_bias; // @[Conv.scala 61:37]
  wire [17:0] addtree_0_io_dout; // @[Conv.scala 61:37]
  wire  addtree_1_clock; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_0; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_1; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_2; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_3; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_4; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_5; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_6; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_din_7; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_bias; // @[Conv.scala 61:37]
  wire [17:0] addtree_1_io_dout; // @[Conv.scala 61:37]
  conv_win_3_3 conv_33_0 ( // @[Conv.scala 47:40]
    .clock(conv_33_0_clock),
    .io_ifm_win_33_0(conv_33_0_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_0_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_0_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_0_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_0_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_0_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_0_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_0_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_0_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_0_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_0_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_0_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_0_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_0_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_0_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_0_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_0_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_0_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_0_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_0_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_0_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_0_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_0_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_0_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_0_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_0_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_0_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_0_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_0_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_1 ( // @[Conv.scala 47:40]
    .clock(conv_33_1_clock),
    .io_ifm_win_33_0(conv_33_1_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_1_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_1_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_1_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_1_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_1_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_1_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_1_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_1_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_1_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_1_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_1_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_1_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_1_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_1_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_1_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_1_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_1_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_1_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_1_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_1_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_1_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_1_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_1_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_1_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_1_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_1_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_1_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_1_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_2 ( // @[Conv.scala 47:40]
    .clock(conv_33_2_clock),
    .io_ifm_win_33_0(conv_33_2_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_2_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_2_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_2_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_2_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_2_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_2_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_2_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_2_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_2_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_2_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_2_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_2_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_2_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_2_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_2_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_2_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_2_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_2_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_2_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_2_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_2_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_2_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_2_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_2_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_2_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_2_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_2_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_2_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_3 ( // @[Conv.scala 47:40]
    .clock(conv_33_3_clock),
    .io_ifm_win_33_0(conv_33_3_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_3_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_3_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_3_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_3_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_3_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_3_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_3_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_3_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_3_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_3_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_3_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_3_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_3_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_3_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_3_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_3_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_3_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_3_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_3_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_3_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_3_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_3_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_3_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_3_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_3_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_3_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_3_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_3_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_4 ( // @[Conv.scala 47:40]
    .clock(conv_33_4_clock),
    .io_ifm_win_33_0(conv_33_4_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_4_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_4_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_4_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_4_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_4_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_4_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_4_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_4_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_4_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_4_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_4_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_4_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_4_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_4_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_4_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_4_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_4_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_4_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_4_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_4_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_4_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_4_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_4_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_4_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_4_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_4_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_4_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_4_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_5 ( // @[Conv.scala 47:40]
    .clock(conv_33_5_clock),
    .io_ifm_win_33_0(conv_33_5_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_5_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_5_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_5_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_5_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_5_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_5_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_5_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_5_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_5_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_5_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_5_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_5_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_5_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_5_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_5_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_5_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_5_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_5_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_5_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_5_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_5_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_5_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_5_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_5_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_5_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_5_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_5_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_5_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_6 ( // @[Conv.scala 47:40]
    .clock(conv_33_6_clock),
    .io_ifm_win_33_0(conv_33_6_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_6_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_6_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_6_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_6_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_6_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_6_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_6_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_6_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_6_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_6_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_6_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_6_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_6_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_6_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_6_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_6_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_6_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_6_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_6_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_6_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_6_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_6_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_6_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_6_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_6_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_6_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_6_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_6_io_o_conv_ch2)
  );
  conv_win_3_3 conv_33_7 ( // @[Conv.scala 47:40]
    .clock(conv_33_7_clock),
    .io_ifm_win_33_0(conv_33_7_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_33_7_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_33_7_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_33_7_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_33_7_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_33_7_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_33_7_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_33_7_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_33_7_io_ifm_win_33_8),
    .io_weight_win_33_ch1_0(conv_33_7_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_33_7_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_33_7_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_33_7_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_33_7_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_33_7_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_33_7_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_33_7_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_33_7_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch2_0(conv_33_7_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_33_7_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_33_7_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_33_7_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_33_7_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_33_7_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_33_7_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_33_7_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_33_7_io_weight_win_33_ch2_8),
    .io_o_conv_ch1(conv_33_7_io_o_conv_ch1),
    .io_o_conv_ch2(conv_33_7_io_o_conv_ch2)
  );
  addtree_int18_3_3 addtree_0 ( // @[Conv.scala 61:37]
    .clock(addtree_0_clock),
    .io_din_0(addtree_0_io_din_0),
    .io_din_1(addtree_0_io_din_1),
    .io_din_2(addtree_0_io_din_2),
    .io_din_3(addtree_0_io_din_3),
    .io_din_4(addtree_0_io_din_4),
    .io_din_5(addtree_0_io_din_5),
    .io_din_6(addtree_0_io_din_6),
    .io_din_7(addtree_0_io_din_7),
    .io_bias(addtree_0_io_bias),
    .io_dout(addtree_0_io_dout)
  );
  addtree_int18_3_3 addtree_1 ( // @[Conv.scala 61:37]
    .clock(addtree_1_clock),
    .io_din_0(addtree_1_io_din_0),
    .io_din_1(addtree_1_io_din_1),
    .io_din_2(addtree_1_io_din_2),
    .io_din_3(addtree_1_io_din_3),
    .io_din_4(addtree_1_io_din_4),
    .io_din_5(addtree_1_io_din_5),
    .io_din_6(addtree_1_io_din_6),
    .io_din_7(addtree_1_io_din_7),
    .io_bias(addtree_1_io_bias),
    .io_dout(addtree_1_io_dout)
  );
  assign io_o_conv_ch1 = addtree_0_io_dout; // @[Conv.scala 68:19]
  assign io_o_conv_ch2 = addtree_1_io_dout; // @[Conv.scala 69:19]
  assign conv_33_0_clock = clock;
  assign conv_33_0_io_ifm_win_33_0 = io_ifm_win_33_0; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_1 = io_ifm_win_33_1; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_2 = io_ifm_win_33_2; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_3 = io_ifm_win_33_3; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_4 = io_ifm_win_33_4; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_5 = io_ifm_win_33_5; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_6 = io_ifm_win_33_6; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_7 = io_ifm_win_33_7; // @[Conv.scala 50:41]
  assign conv_33_0_io_ifm_win_33_8 = io_ifm_win_33_8; // @[Conv.scala 50:41]
  assign conv_33_0_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_0; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_1; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_2; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_3; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_4; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_5; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_6; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_7; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_8; // @[Conv.scala 51:48]
  assign conv_33_0_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_0; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_1; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_2; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_3; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_4; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_5; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_6; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_7; // @[Conv.scala 52:48]
  assign conv_33_0_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_8; // @[Conv.scala 52:48]
  assign conv_33_1_clock = clock;
  assign conv_33_1_io_ifm_win_33_0 = io_ifm_win_33_9; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_1 = io_ifm_win_33_10; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_2 = io_ifm_win_33_11; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_3 = io_ifm_win_33_12; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_4 = io_ifm_win_33_13; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_5 = io_ifm_win_33_14; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_6 = io_ifm_win_33_15; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_7 = io_ifm_win_33_16; // @[Conv.scala 50:41]
  assign conv_33_1_io_ifm_win_33_8 = io_ifm_win_33_17; // @[Conv.scala 50:41]
  assign conv_33_1_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_9; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_10; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_11; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_12; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_13; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_14; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_15; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_16; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_17; // @[Conv.scala 51:48]
  assign conv_33_1_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_9; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_10; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_11; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_12; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_13; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_14; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_15; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_16; // @[Conv.scala 52:48]
  assign conv_33_1_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_17; // @[Conv.scala 52:48]
  assign conv_33_2_clock = clock;
  assign conv_33_2_io_ifm_win_33_0 = io_ifm_win_33_18; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_1 = io_ifm_win_33_19; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_2 = io_ifm_win_33_20; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_3 = io_ifm_win_33_21; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_4 = io_ifm_win_33_22; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_5 = io_ifm_win_33_23; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_6 = io_ifm_win_33_24; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_7 = io_ifm_win_33_25; // @[Conv.scala 50:41]
  assign conv_33_2_io_ifm_win_33_8 = io_ifm_win_33_26; // @[Conv.scala 50:41]
  assign conv_33_2_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_18; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_19; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_20; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_21; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_22; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_23; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_24; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_25; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_26; // @[Conv.scala 51:48]
  assign conv_33_2_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_18; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_19; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_20; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_21; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_22; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_23; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_24; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_25; // @[Conv.scala 52:48]
  assign conv_33_2_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_26; // @[Conv.scala 52:48]
  assign conv_33_3_clock = clock;
  assign conv_33_3_io_ifm_win_33_0 = io_ifm_win_33_27; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_1 = io_ifm_win_33_28; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_2 = io_ifm_win_33_29; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_3 = io_ifm_win_33_30; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_4 = io_ifm_win_33_31; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_5 = io_ifm_win_33_32; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_6 = io_ifm_win_33_33; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_7 = io_ifm_win_33_34; // @[Conv.scala 50:41]
  assign conv_33_3_io_ifm_win_33_8 = io_ifm_win_33_35; // @[Conv.scala 50:41]
  assign conv_33_3_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_27; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_28; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_29; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_30; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_31; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_32; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_33; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_34; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_35; // @[Conv.scala 51:48]
  assign conv_33_3_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_27; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_28; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_29; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_30; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_31; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_32; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_33; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_34; // @[Conv.scala 52:48]
  assign conv_33_3_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_35; // @[Conv.scala 52:48]
  assign conv_33_4_clock = clock;
  assign conv_33_4_io_ifm_win_33_0 = io_ifm_win_33_36; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_1 = io_ifm_win_33_37; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_2 = io_ifm_win_33_38; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_3 = io_ifm_win_33_39; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_4 = io_ifm_win_33_40; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_5 = io_ifm_win_33_41; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_6 = io_ifm_win_33_42; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_7 = io_ifm_win_33_43; // @[Conv.scala 50:41]
  assign conv_33_4_io_ifm_win_33_8 = io_ifm_win_33_44; // @[Conv.scala 50:41]
  assign conv_33_4_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_36; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_37; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_38; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_39; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_40; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_41; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_42; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_43; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_44; // @[Conv.scala 51:48]
  assign conv_33_4_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_36; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_37; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_38; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_39; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_40; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_41; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_42; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_43; // @[Conv.scala 52:48]
  assign conv_33_4_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_44; // @[Conv.scala 52:48]
  assign conv_33_5_clock = clock;
  assign conv_33_5_io_ifm_win_33_0 = io_ifm_win_33_45; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_1 = io_ifm_win_33_46; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_2 = io_ifm_win_33_47; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_3 = io_ifm_win_33_48; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_4 = io_ifm_win_33_49; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_5 = io_ifm_win_33_50; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_6 = io_ifm_win_33_51; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_7 = io_ifm_win_33_52; // @[Conv.scala 50:41]
  assign conv_33_5_io_ifm_win_33_8 = io_ifm_win_33_53; // @[Conv.scala 50:41]
  assign conv_33_5_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_45; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_46; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_47; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_48; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_49; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_50; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_51; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_52; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_53; // @[Conv.scala 51:48]
  assign conv_33_5_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_45; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_46; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_47; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_48; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_49; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_50; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_51; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_52; // @[Conv.scala 52:48]
  assign conv_33_5_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_53; // @[Conv.scala 52:48]
  assign conv_33_6_clock = clock;
  assign conv_33_6_io_ifm_win_33_0 = io_ifm_win_33_54; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_1 = io_ifm_win_33_55; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_2 = io_ifm_win_33_56; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_3 = io_ifm_win_33_57; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_4 = io_ifm_win_33_58; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_5 = io_ifm_win_33_59; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_6 = io_ifm_win_33_60; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_7 = io_ifm_win_33_61; // @[Conv.scala 50:41]
  assign conv_33_6_io_ifm_win_33_8 = io_ifm_win_33_62; // @[Conv.scala 50:41]
  assign conv_33_6_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_54; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_55; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_56; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_57; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_58; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_59; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_60; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_61; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_62; // @[Conv.scala 51:48]
  assign conv_33_6_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_54; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_55; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_56; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_57; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_58; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_59; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_60; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_61; // @[Conv.scala 52:48]
  assign conv_33_6_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_62; // @[Conv.scala 52:48]
  assign conv_33_7_clock = clock;
  assign conv_33_7_io_ifm_win_33_0 = io_ifm_win_33_63; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_1 = io_ifm_win_33_64; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_2 = io_ifm_win_33_65; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_3 = io_ifm_win_33_66; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_4 = io_ifm_win_33_67; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_5 = io_ifm_win_33_68; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_6 = io_ifm_win_33_69; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_7 = io_ifm_win_33_70; // @[Conv.scala 50:41]
  assign conv_33_7_io_ifm_win_33_8 = io_ifm_win_33_71; // @[Conv.scala 50:41]
  assign conv_33_7_io_weight_win_33_ch1_0 = io_weight_win_33_ch1_63; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_1 = io_weight_win_33_ch1_64; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_2 = io_weight_win_33_ch1_65; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_3 = io_weight_win_33_ch1_66; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_4 = io_weight_win_33_ch1_67; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_5 = io_weight_win_33_ch1_68; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_6 = io_weight_win_33_ch1_69; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_7 = io_weight_win_33_ch1_70; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch1_8 = io_weight_win_33_ch1_71; // @[Conv.scala 51:48]
  assign conv_33_7_io_weight_win_33_ch2_0 = io_weight_win_33_ch2_63; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_1 = io_weight_win_33_ch2_64; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_2 = io_weight_win_33_ch2_65; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_3 = io_weight_win_33_ch2_66; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_4 = io_weight_win_33_ch2_67; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_5 = io_weight_win_33_ch2_68; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_6 = io_weight_win_33_ch2_69; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_7 = io_weight_win_33_ch2_70; // @[Conv.scala 52:48]
  assign conv_33_7_io_weight_win_33_ch2_8 = io_weight_win_33_ch2_71; // @[Conv.scala 52:48]
  assign addtree_0_clock = clock;
  assign addtree_0_io_din_0 = conv_33_0_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_1 = conv_33_1_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_2 = conv_33_2_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_3 = conv_33_3_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_4 = conv_33_4_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_5 = conv_33_5_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_6 = conv_33_6_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_din_7 = conv_33_7_io_o_conv_ch1; // @[Conv.scala 45:19 54:16]
  assign addtree_0_io_bias = io_bias_valid ? io_bias1 : 18'h0; // @[Conv.scala 58:23]
  assign addtree_1_clock = clock;
  assign addtree_1_io_din_0 = conv_33_0_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_1 = conv_33_1_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_2 = conv_33_2_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_3 = conv_33_3_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_4 = conv_33_4_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_5 = conv_33_5_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_6 = conv_33_6_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_din_7 = conv_33_7_io_o_conv_ch2; // @[Conv.scala 46:19 55:16]
  assign addtree_1_io_bias = io_bias_valid ? io_bias2 : 18'h0; // @[Conv.scala 59:23]
endmodule
module Conv(
  input         clock,
  input  [7:0]  io_ifm_win_33_0,
  input  [7:0]  io_ifm_win_33_1,
  input  [7:0]  io_ifm_win_33_2,
  input  [7:0]  io_ifm_win_33_3,
  input  [7:0]  io_ifm_win_33_4,
  input  [7:0]  io_ifm_win_33_5,
  input  [7:0]  io_ifm_win_33_6,
  input  [7:0]  io_ifm_win_33_7,
  input  [7:0]  io_ifm_win_33_8,
  input  [7:0]  io_ifm_win_33_9,
  input  [7:0]  io_ifm_win_33_10,
  input  [7:0]  io_ifm_win_33_11,
  input  [7:0]  io_ifm_win_33_12,
  input  [7:0]  io_ifm_win_33_13,
  input  [7:0]  io_ifm_win_33_14,
  input  [7:0]  io_ifm_win_33_15,
  input  [7:0]  io_ifm_win_33_16,
  input  [7:0]  io_ifm_win_33_17,
  input  [7:0]  io_ifm_win_33_18,
  input  [7:0]  io_ifm_win_33_19,
  input  [7:0]  io_ifm_win_33_20,
  input  [7:0]  io_ifm_win_33_21,
  input  [7:0]  io_ifm_win_33_22,
  input  [7:0]  io_ifm_win_33_23,
  input  [7:0]  io_ifm_win_33_24,
  input  [7:0]  io_ifm_win_33_25,
  input  [7:0]  io_ifm_win_33_26,
  input  [7:0]  io_ifm_win_33_27,
  input  [7:0]  io_ifm_win_33_28,
  input  [7:0]  io_ifm_win_33_29,
  input  [7:0]  io_ifm_win_33_30,
  input  [7:0]  io_ifm_win_33_31,
  input  [7:0]  io_ifm_win_33_32,
  input  [7:0]  io_ifm_win_33_33,
  input  [7:0]  io_ifm_win_33_34,
  input  [7:0]  io_ifm_win_33_35,
  input  [7:0]  io_ifm_win_33_36,
  input  [7:0]  io_ifm_win_33_37,
  input  [7:0]  io_ifm_win_33_38,
  input  [7:0]  io_ifm_win_33_39,
  input  [7:0]  io_ifm_win_33_40,
  input  [7:0]  io_ifm_win_33_41,
  input  [7:0]  io_ifm_win_33_42,
  input  [7:0]  io_ifm_win_33_43,
  input  [7:0]  io_ifm_win_33_44,
  input  [7:0]  io_ifm_win_33_45,
  input  [7:0]  io_ifm_win_33_46,
  input  [7:0]  io_ifm_win_33_47,
  input  [7:0]  io_ifm_win_33_48,
  input  [7:0]  io_ifm_win_33_49,
  input  [7:0]  io_ifm_win_33_50,
  input  [7:0]  io_ifm_win_33_51,
  input  [7:0]  io_ifm_win_33_52,
  input  [7:0]  io_ifm_win_33_53,
  input  [7:0]  io_ifm_win_33_54,
  input  [7:0]  io_ifm_win_33_55,
  input  [7:0]  io_ifm_win_33_56,
  input  [7:0]  io_ifm_win_33_57,
  input  [7:0]  io_ifm_win_33_58,
  input  [7:0]  io_ifm_win_33_59,
  input  [7:0]  io_ifm_win_33_60,
  input  [7:0]  io_ifm_win_33_61,
  input  [7:0]  io_ifm_win_33_62,
  input  [7:0]  io_ifm_win_33_63,
  input  [7:0]  io_ifm_win_33_64,
  input  [7:0]  io_ifm_win_33_65,
  input  [7:0]  io_ifm_win_33_66,
  input  [7:0]  io_ifm_win_33_67,
  input  [7:0]  io_ifm_win_33_68,
  input  [7:0]  io_ifm_win_33_69,
  input  [7:0]  io_ifm_win_33_70,
  input  [7:0]  io_ifm_win_33_71,
  input  [7:0]  io_weight_win_33_0,
  input  [7:0]  io_weight_win_33_1,
  input  [7:0]  io_weight_win_33_2,
  input  [7:0]  io_weight_win_33_3,
  input  [7:0]  io_weight_win_33_4,
  input  [7:0]  io_weight_win_33_5,
  input  [7:0]  io_weight_win_33_6,
  input  [7:0]  io_weight_win_33_7,
  input  [7:0]  io_weight_win_33_8,
  input  [7:0]  io_weight_win_33_9,
  input  [7:0]  io_weight_win_33_10,
  input  [7:0]  io_weight_win_33_11,
  input  [7:0]  io_weight_win_33_12,
  input  [7:0]  io_weight_win_33_13,
  input  [7:0]  io_weight_win_33_14,
  input  [7:0]  io_weight_win_33_15,
  input  [7:0]  io_weight_win_33_16,
  input  [7:0]  io_weight_win_33_17,
  input  [7:0]  io_weight_win_33_18,
  input  [7:0]  io_weight_win_33_19,
  input  [7:0]  io_weight_win_33_20,
  input  [7:0]  io_weight_win_33_21,
  input  [7:0]  io_weight_win_33_22,
  input  [7:0]  io_weight_win_33_23,
  input  [7:0]  io_weight_win_33_24,
  input  [7:0]  io_weight_win_33_25,
  input  [7:0]  io_weight_win_33_26,
  input  [7:0]  io_weight_win_33_27,
  input  [7:0]  io_weight_win_33_28,
  input  [7:0]  io_weight_win_33_29,
  input  [7:0]  io_weight_win_33_30,
  input  [7:0]  io_weight_win_33_31,
  input  [7:0]  io_weight_win_33_32,
  input  [7:0]  io_weight_win_33_33,
  input  [7:0]  io_weight_win_33_34,
  input  [7:0]  io_weight_win_33_35,
  input  [7:0]  io_weight_win_33_36,
  input  [7:0]  io_weight_win_33_37,
  input  [7:0]  io_weight_win_33_38,
  input  [7:0]  io_weight_win_33_39,
  input  [7:0]  io_weight_win_33_40,
  input  [7:0]  io_weight_win_33_41,
  input  [7:0]  io_weight_win_33_42,
  input  [7:0]  io_weight_win_33_43,
  input  [7:0]  io_weight_win_33_44,
  input  [7:0]  io_weight_win_33_45,
  input  [7:0]  io_weight_win_33_46,
  input  [7:0]  io_weight_win_33_47,
  input  [7:0]  io_weight_win_33_48,
  input  [7:0]  io_weight_win_33_49,
  input  [7:0]  io_weight_win_33_50,
  input  [7:0]  io_weight_win_33_51,
  input  [7:0]  io_weight_win_33_52,
  input  [7:0]  io_weight_win_33_53,
  input  [7:0]  io_weight_win_33_54,
  input  [7:0]  io_weight_win_33_55,
  input  [7:0]  io_weight_win_33_56,
  input  [7:0]  io_weight_win_33_57,
  input  [7:0]  io_weight_win_33_58,
  input  [7:0]  io_weight_win_33_59,
  input  [7:0]  io_weight_win_33_60,
  input  [7:0]  io_weight_win_33_61,
  input  [7:0]  io_weight_win_33_62,
  input  [7:0]  io_weight_win_33_63,
  input  [7:0]  io_weight_win_33_64,
  input  [7:0]  io_weight_win_33_65,
  input  [7:0]  io_weight_win_33_66,
  input  [7:0]  io_weight_win_33_67,
  input  [7:0]  io_weight_win_33_68,
  input  [7:0]  io_weight_win_33_69,
  input  [7:0]  io_weight_win_33_70,
  input  [7:0]  io_weight_win_33_71,
  input  [7:0]  io_weight_win_33_72,
  input  [7:0]  io_weight_win_33_73,
  input  [7:0]  io_weight_win_33_74,
  input  [7:0]  io_weight_win_33_75,
  input  [7:0]  io_weight_win_33_76,
  input  [7:0]  io_weight_win_33_77,
  input  [7:0]  io_weight_win_33_78,
  input  [7:0]  io_weight_win_33_79,
  input  [7:0]  io_weight_win_33_80,
  input  [7:0]  io_weight_win_33_81,
  input  [7:0]  io_weight_win_33_82,
  input  [7:0]  io_weight_win_33_83,
  input  [7:0]  io_weight_win_33_84,
  input  [7:0]  io_weight_win_33_85,
  input  [7:0]  io_weight_win_33_86,
  input  [7:0]  io_weight_win_33_87,
  input  [7:0]  io_weight_win_33_88,
  input  [7:0]  io_weight_win_33_89,
  input  [7:0]  io_weight_win_33_90,
  input  [7:0]  io_weight_win_33_91,
  input  [7:0]  io_weight_win_33_92,
  input  [7:0]  io_weight_win_33_93,
  input  [7:0]  io_weight_win_33_94,
  input  [7:0]  io_weight_win_33_95,
  input  [7:0]  io_weight_win_33_96,
  input  [7:0]  io_weight_win_33_97,
  input  [7:0]  io_weight_win_33_98,
  input  [7:0]  io_weight_win_33_99,
  input  [7:0]  io_weight_win_33_100,
  input  [7:0]  io_weight_win_33_101,
  input  [7:0]  io_weight_win_33_102,
  input  [7:0]  io_weight_win_33_103,
  input  [7:0]  io_weight_win_33_104,
  input  [7:0]  io_weight_win_33_105,
  input  [7:0]  io_weight_win_33_106,
  input  [7:0]  io_weight_win_33_107,
  input  [7:0]  io_weight_win_33_108,
  input  [7:0]  io_weight_win_33_109,
  input  [7:0]  io_weight_win_33_110,
  input  [7:0]  io_weight_win_33_111,
  input  [7:0]  io_weight_win_33_112,
  input  [7:0]  io_weight_win_33_113,
  input  [7:0]  io_weight_win_33_114,
  input  [7:0]  io_weight_win_33_115,
  input  [7:0]  io_weight_win_33_116,
  input  [7:0]  io_weight_win_33_117,
  input  [7:0]  io_weight_win_33_118,
  input  [7:0]  io_weight_win_33_119,
  input  [7:0]  io_weight_win_33_120,
  input  [7:0]  io_weight_win_33_121,
  input  [7:0]  io_weight_win_33_122,
  input  [7:0]  io_weight_win_33_123,
  input  [7:0]  io_weight_win_33_124,
  input  [7:0]  io_weight_win_33_125,
  input  [7:0]  io_weight_win_33_126,
  input  [7:0]  io_weight_win_33_127,
  input  [7:0]  io_weight_win_33_128,
  input  [7:0]  io_weight_win_33_129,
  input  [7:0]  io_weight_win_33_130,
  input  [7:0]  io_weight_win_33_131,
  input  [7:0]  io_weight_win_33_132,
  input  [7:0]  io_weight_win_33_133,
  input  [7:0]  io_weight_win_33_134,
  input  [7:0]  io_weight_win_33_135,
  input  [7:0]  io_weight_win_33_136,
  input  [7:0]  io_weight_win_33_137,
  input  [7:0]  io_weight_win_33_138,
  input  [7:0]  io_weight_win_33_139,
  input  [7:0]  io_weight_win_33_140,
  input  [7:0]  io_weight_win_33_141,
  input  [7:0]  io_weight_win_33_142,
  input  [7:0]  io_weight_win_33_143,
  input  [7:0]  io_weight_win_33_144,
  input  [7:0]  io_weight_win_33_145,
  input  [7:0]  io_weight_win_33_146,
  input  [7:0]  io_weight_win_33_147,
  input  [7:0]  io_weight_win_33_148,
  input  [7:0]  io_weight_win_33_149,
  input  [7:0]  io_weight_win_33_150,
  input  [7:0]  io_weight_win_33_151,
  input  [7:0]  io_weight_win_33_152,
  input  [7:0]  io_weight_win_33_153,
  input  [7:0]  io_weight_win_33_154,
  input  [7:0]  io_weight_win_33_155,
  input  [7:0]  io_weight_win_33_156,
  input  [7:0]  io_weight_win_33_157,
  input  [7:0]  io_weight_win_33_158,
  input  [7:0]  io_weight_win_33_159,
  input  [7:0]  io_weight_win_33_160,
  input  [7:0]  io_weight_win_33_161,
  input  [7:0]  io_weight_win_33_162,
  input  [7:0]  io_weight_win_33_163,
  input  [7:0]  io_weight_win_33_164,
  input  [7:0]  io_weight_win_33_165,
  input  [7:0]  io_weight_win_33_166,
  input  [7:0]  io_weight_win_33_167,
  input  [7:0]  io_weight_win_33_168,
  input  [7:0]  io_weight_win_33_169,
  input  [7:0]  io_weight_win_33_170,
  input  [7:0]  io_weight_win_33_171,
  input  [7:0]  io_weight_win_33_172,
  input  [7:0]  io_weight_win_33_173,
  input  [7:0]  io_weight_win_33_174,
  input  [7:0]  io_weight_win_33_175,
  input  [7:0]  io_weight_win_33_176,
  input  [7:0]  io_weight_win_33_177,
  input  [7:0]  io_weight_win_33_178,
  input  [7:0]  io_weight_win_33_179,
  input  [7:0]  io_weight_win_33_180,
  input  [7:0]  io_weight_win_33_181,
  input  [7:0]  io_weight_win_33_182,
  input  [7:0]  io_weight_win_33_183,
  input  [7:0]  io_weight_win_33_184,
  input  [7:0]  io_weight_win_33_185,
  input  [7:0]  io_weight_win_33_186,
  input  [7:0]  io_weight_win_33_187,
  input  [7:0]  io_weight_win_33_188,
  input  [7:0]  io_weight_win_33_189,
  input  [7:0]  io_weight_win_33_190,
  input  [7:0]  io_weight_win_33_191,
  input  [7:0]  io_weight_win_33_192,
  input  [7:0]  io_weight_win_33_193,
  input  [7:0]  io_weight_win_33_194,
  input  [7:0]  io_weight_win_33_195,
  input  [7:0]  io_weight_win_33_196,
  input  [7:0]  io_weight_win_33_197,
  input  [7:0]  io_weight_win_33_198,
  input  [7:0]  io_weight_win_33_199,
  input  [7:0]  io_weight_win_33_200,
  input  [7:0]  io_weight_win_33_201,
  input  [7:0]  io_weight_win_33_202,
  input  [7:0]  io_weight_win_33_203,
  input  [7:0]  io_weight_win_33_204,
  input  [7:0]  io_weight_win_33_205,
  input  [7:0]  io_weight_win_33_206,
  input  [7:0]  io_weight_win_33_207,
  input  [7:0]  io_weight_win_33_208,
  input  [7:0]  io_weight_win_33_209,
  input  [7:0]  io_weight_win_33_210,
  input  [7:0]  io_weight_win_33_211,
  input  [7:0]  io_weight_win_33_212,
  input  [7:0]  io_weight_win_33_213,
  input  [7:0]  io_weight_win_33_214,
  input  [7:0]  io_weight_win_33_215,
  input  [7:0]  io_weight_win_33_216,
  input  [7:0]  io_weight_win_33_217,
  input  [7:0]  io_weight_win_33_218,
  input  [7:0]  io_weight_win_33_219,
  input  [7:0]  io_weight_win_33_220,
  input  [7:0]  io_weight_win_33_221,
  input  [7:0]  io_weight_win_33_222,
  input  [7:0]  io_weight_win_33_223,
  input  [7:0]  io_weight_win_33_224,
  input  [7:0]  io_weight_win_33_225,
  input  [7:0]  io_weight_win_33_226,
  input  [7:0]  io_weight_win_33_227,
  input  [7:0]  io_weight_win_33_228,
  input  [7:0]  io_weight_win_33_229,
  input  [7:0]  io_weight_win_33_230,
  input  [7:0]  io_weight_win_33_231,
  input  [7:0]  io_weight_win_33_232,
  input  [7:0]  io_weight_win_33_233,
  input  [7:0]  io_weight_win_33_234,
  input  [7:0]  io_weight_win_33_235,
  input  [7:0]  io_weight_win_33_236,
  input  [7:0]  io_weight_win_33_237,
  input  [7:0]  io_weight_win_33_238,
  input  [7:0]  io_weight_win_33_239,
  input  [7:0]  io_weight_win_33_240,
  input  [7:0]  io_weight_win_33_241,
  input  [7:0]  io_weight_win_33_242,
  input  [7:0]  io_weight_win_33_243,
  input  [7:0]  io_weight_win_33_244,
  input  [7:0]  io_weight_win_33_245,
  input  [7:0]  io_weight_win_33_246,
  input  [7:0]  io_weight_win_33_247,
  input  [7:0]  io_weight_win_33_248,
  input  [7:0]  io_weight_win_33_249,
  input  [7:0]  io_weight_win_33_250,
  input  [7:0]  io_weight_win_33_251,
  input  [7:0]  io_weight_win_33_252,
  input  [7:0]  io_weight_win_33_253,
  input  [7:0]  io_weight_win_33_254,
  input  [7:0]  io_weight_win_33_255,
  input  [7:0]  io_weight_win_33_256,
  input  [7:0]  io_weight_win_33_257,
  input  [7:0]  io_weight_win_33_258,
  input  [7:0]  io_weight_win_33_259,
  input  [7:0]  io_weight_win_33_260,
  input  [7:0]  io_weight_win_33_261,
  input  [7:0]  io_weight_win_33_262,
  input  [7:0]  io_weight_win_33_263,
  input  [7:0]  io_weight_win_33_264,
  input  [7:0]  io_weight_win_33_265,
  input  [7:0]  io_weight_win_33_266,
  input  [7:0]  io_weight_win_33_267,
  input  [7:0]  io_weight_win_33_268,
  input  [7:0]  io_weight_win_33_269,
  input  [7:0]  io_weight_win_33_270,
  input  [7:0]  io_weight_win_33_271,
  input  [7:0]  io_weight_win_33_272,
  input  [7:0]  io_weight_win_33_273,
  input  [7:0]  io_weight_win_33_274,
  input  [7:0]  io_weight_win_33_275,
  input  [7:0]  io_weight_win_33_276,
  input  [7:0]  io_weight_win_33_277,
  input  [7:0]  io_weight_win_33_278,
  input  [7:0]  io_weight_win_33_279,
  input  [7:0]  io_weight_win_33_280,
  input  [7:0]  io_weight_win_33_281,
  input  [7:0]  io_weight_win_33_282,
  input  [7:0]  io_weight_win_33_283,
  input  [7:0]  io_weight_win_33_284,
  input  [7:0]  io_weight_win_33_285,
  input  [7:0]  io_weight_win_33_286,
  input  [7:0]  io_weight_win_33_287,
  input  [7:0]  io_weight_win_33_288,
  input  [7:0]  io_weight_win_33_289,
  input  [7:0]  io_weight_win_33_290,
  input  [7:0]  io_weight_win_33_291,
  input  [7:0]  io_weight_win_33_292,
  input  [7:0]  io_weight_win_33_293,
  input  [7:0]  io_weight_win_33_294,
  input  [7:0]  io_weight_win_33_295,
  input  [7:0]  io_weight_win_33_296,
  input  [7:0]  io_weight_win_33_297,
  input  [7:0]  io_weight_win_33_298,
  input  [7:0]  io_weight_win_33_299,
  input  [7:0]  io_weight_win_33_300,
  input  [7:0]  io_weight_win_33_301,
  input  [7:0]  io_weight_win_33_302,
  input  [7:0]  io_weight_win_33_303,
  input  [7:0]  io_weight_win_33_304,
  input  [7:0]  io_weight_win_33_305,
  input  [7:0]  io_weight_win_33_306,
  input  [7:0]  io_weight_win_33_307,
  input  [7:0]  io_weight_win_33_308,
  input  [7:0]  io_weight_win_33_309,
  input  [7:0]  io_weight_win_33_310,
  input  [7:0]  io_weight_win_33_311,
  input  [7:0]  io_weight_win_33_312,
  input  [7:0]  io_weight_win_33_313,
  input  [7:0]  io_weight_win_33_314,
  input  [7:0]  io_weight_win_33_315,
  input  [7:0]  io_weight_win_33_316,
  input  [7:0]  io_weight_win_33_317,
  input  [7:0]  io_weight_win_33_318,
  input  [7:0]  io_weight_win_33_319,
  input  [7:0]  io_weight_win_33_320,
  input  [7:0]  io_weight_win_33_321,
  input  [7:0]  io_weight_win_33_322,
  input  [7:0]  io_weight_win_33_323,
  input  [7:0]  io_weight_win_33_324,
  input  [7:0]  io_weight_win_33_325,
  input  [7:0]  io_weight_win_33_326,
  input  [7:0]  io_weight_win_33_327,
  input  [7:0]  io_weight_win_33_328,
  input  [7:0]  io_weight_win_33_329,
  input  [7:0]  io_weight_win_33_330,
  input  [7:0]  io_weight_win_33_331,
  input  [7:0]  io_weight_win_33_332,
  input  [7:0]  io_weight_win_33_333,
  input  [7:0]  io_weight_win_33_334,
  input  [7:0]  io_weight_win_33_335,
  input  [7:0]  io_weight_win_33_336,
  input  [7:0]  io_weight_win_33_337,
  input  [7:0]  io_weight_win_33_338,
  input  [7:0]  io_weight_win_33_339,
  input  [7:0]  io_weight_win_33_340,
  input  [7:0]  io_weight_win_33_341,
  input  [7:0]  io_weight_win_33_342,
  input  [7:0]  io_weight_win_33_343,
  input  [7:0]  io_weight_win_33_344,
  input  [7:0]  io_weight_win_33_345,
  input  [7:0]  io_weight_win_33_346,
  input  [7:0]  io_weight_win_33_347,
  input  [7:0]  io_weight_win_33_348,
  input  [7:0]  io_weight_win_33_349,
  input  [7:0]  io_weight_win_33_350,
  input  [7:0]  io_weight_win_33_351,
  input  [7:0]  io_weight_win_33_352,
  input  [7:0]  io_weight_win_33_353,
  input  [7:0]  io_weight_win_33_354,
  input  [7:0]  io_weight_win_33_355,
  input  [7:0]  io_weight_win_33_356,
  input  [7:0]  io_weight_win_33_357,
  input  [7:0]  io_weight_win_33_358,
  input  [7:0]  io_weight_win_33_359,
  input  [7:0]  io_weight_win_33_360,
  input  [7:0]  io_weight_win_33_361,
  input  [7:0]  io_weight_win_33_362,
  input  [7:0]  io_weight_win_33_363,
  input  [7:0]  io_weight_win_33_364,
  input  [7:0]  io_weight_win_33_365,
  input  [7:0]  io_weight_win_33_366,
  input  [7:0]  io_weight_win_33_367,
  input  [7:0]  io_weight_win_33_368,
  input  [7:0]  io_weight_win_33_369,
  input  [7:0]  io_weight_win_33_370,
  input  [7:0]  io_weight_win_33_371,
  input  [7:0]  io_weight_win_33_372,
  input  [7:0]  io_weight_win_33_373,
  input  [7:0]  io_weight_win_33_374,
  input  [7:0]  io_weight_win_33_375,
  input  [7:0]  io_weight_win_33_376,
  input  [7:0]  io_weight_win_33_377,
  input  [7:0]  io_weight_win_33_378,
  input  [7:0]  io_weight_win_33_379,
  input  [7:0]  io_weight_win_33_380,
  input  [7:0]  io_weight_win_33_381,
  input  [7:0]  io_weight_win_33_382,
  input  [7:0]  io_weight_win_33_383,
  input  [7:0]  io_weight_win_33_384,
  input  [7:0]  io_weight_win_33_385,
  input  [7:0]  io_weight_win_33_386,
  input  [7:0]  io_weight_win_33_387,
  input  [7:0]  io_weight_win_33_388,
  input  [7:0]  io_weight_win_33_389,
  input  [7:0]  io_weight_win_33_390,
  input  [7:0]  io_weight_win_33_391,
  input  [7:0]  io_weight_win_33_392,
  input  [7:0]  io_weight_win_33_393,
  input  [7:0]  io_weight_win_33_394,
  input  [7:0]  io_weight_win_33_395,
  input  [7:0]  io_weight_win_33_396,
  input  [7:0]  io_weight_win_33_397,
  input  [7:0]  io_weight_win_33_398,
  input  [7:0]  io_weight_win_33_399,
  input  [7:0]  io_weight_win_33_400,
  input  [7:0]  io_weight_win_33_401,
  input  [7:0]  io_weight_win_33_402,
  input  [7:0]  io_weight_win_33_403,
  input  [7:0]  io_weight_win_33_404,
  input  [7:0]  io_weight_win_33_405,
  input  [7:0]  io_weight_win_33_406,
  input  [7:0]  io_weight_win_33_407,
  input  [7:0]  io_weight_win_33_408,
  input  [7:0]  io_weight_win_33_409,
  input  [7:0]  io_weight_win_33_410,
  input  [7:0]  io_weight_win_33_411,
  input  [7:0]  io_weight_win_33_412,
  input  [7:0]  io_weight_win_33_413,
  input  [7:0]  io_weight_win_33_414,
  input  [7:0]  io_weight_win_33_415,
  input  [7:0]  io_weight_win_33_416,
  input  [7:0]  io_weight_win_33_417,
  input  [7:0]  io_weight_win_33_418,
  input  [7:0]  io_weight_win_33_419,
  input  [7:0]  io_weight_win_33_420,
  input  [7:0]  io_weight_win_33_421,
  input  [7:0]  io_weight_win_33_422,
  input  [7:0]  io_weight_win_33_423,
  input  [7:0]  io_weight_win_33_424,
  input  [7:0]  io_weight_win_33_425,
  input  [7:0]  io_weight_win_33_426,
  input  [7:0]  io_weight_win_33_427,
  input  [7:0]  io_weight_win_33_428,
  input  [7:0]  io_weight_win_33_429,
  input  [7:0]  io_weight_win_33_430,
  input  [7:0]  io_weight_win_33_431,
  input  [7:0]  io_weight_win_33_432,
  input  [7:0]  io_weight_win_33_433,
  input  [7:0]  io_weight_win_33_434,
  input  [7:0]  io_weight_win_33_435,
  input  [7:0]  io_weight_win_33_436,
  input  [7:0]  io_weight_win_33_437,
  input  [7:0]  io_weight_win_33_438,
  input  [7:0]  io_weight_win_33_439,
  input  [7:0]  io_weight_win_33_440,
  input  [7:0]  io_weight_win_33_441,
  input  [7:0]  io_weight_win_33_442,
  input  [7:0]  io_weight_win_33_443,
  input  [7:0]  io_weight_win_33_444,
  input  [7:0]  io_weight_win_33_445,
  input  [7:0]  io_weight_win_33_446,
  input  [7:0]  io_weight_win_33_447,
  input  [7:0]  io_weight_win_33_448,
  input  [7:0]  io_weight_win_33_449,
  input  [7:0]  io_weight_win_33_450,
  input  [7:0]  io_weight_win_33_451,
  input  [7:0]  io_weight_win_33_452,
  input  [7:0]  io_weight_win_33_453,
  input  [7:0]  io_weight_win_33_454,
  input  [7:0]  io_weight_win_33_455,
  input  [7:0]  io_weight_win_33_456,
  input  [7:0]  io_weight_win_33_457,
  input  [7:0]  io_weight_win_33_458,
  input  [7:0]  io_weight_win_33_459,
  input  [7:0]  io_weight_win_33_460,
  input  [7:0]  io_weight_win_33_461,
  input  [7:0]  io_weight_win_33_462,
  input  [7:0]  io_weight_win_33_463,
  input  [7:0]  io_weight_win_33_464,
  input  [7:0]  io_weight_win_33_465,
  input  [7:0]  io_weight_win_33_466,
  input  [7:0]  io_weight_win_33_467,
  input  [7:0]  io_weight_win_33_468,
  input  [7:0]  io_weight_win_33_469,
  input  [7:0]  io_weight_win_33_470,
  input  [7:0]  io_weight_win_33_471,
  input  [7:0]  io_weight_win_33_472,
  input  [7:0]  io_weight_win_33_473,
  input  [7:0]  io_weight_win_33_474,
  input  [7:0]  io_weight_win_33_475,
  input  [7:0]  io_weight_win_33_476,
  input  [7:0]  io_weight_win_33_477,
  input  [7:0]  io_weight_win_33_478,
  input  [7:0]  io_weight_win_33_479,
  input  [7:0]  io_weight_win_33_480,
  input  [7:0]  io_weight_win_33_481,
  input  [7:0]  io_weight_win_33_482,
  input  [7:0]  io_weight_win_33_483,
  input  [7:0]  io_weight_win_33_484,
  input  [7:0]  io_weight_win_33_485,
  input  [7:0]  io_weight_win_33_486,
  input  [7:0]  io_weight_win_33_487,
  input  [7:0]  io_weight_win_33_488,
  input  [7:0]  io_weight_win_33_489,
  input  [7:0]  io_weight_win_33_490,
  input  [7:0]  io_weight_win_33_491,
  input  [7:0]  io_weight_win_33_492,
  input  [7:0]  io_weight_win_33_493,
  input  [7:0]  io_weight_win_33_494,
  input  [7:0]  io_weight_win_33_495,
  input  [7:0]  io_weight_win_33_496,
  input  [7:0]  io_weight_win_33_497,
  input  [7:0]  io_weight_win_33_498,
  input  [7:0]  io_weight_win_33_499,
  input  [7:0]  io_weight_win_33_500,
  input  [7:0]  io_weight_win_33_501,
  input  [7:0]  io_weight_win_33_502,
  input  [7:0]  io_weight_win_33_503,
  input  [7:0]  io_weight_win_33_504,
  input  [7:0]  io_weight_win_33_505,
  input  [7:0]  io_weight_win_33_506,
  input  [7:0]  io_weight_win_33_507,
  input  [7:0]  io_weight_win_33_508,
  input  [7:0]  io_weight_win_33_509,
  input  [7:0]  io_weight_win_33_510,
  input  [7:0]  io_weight_win_33_511,
  input  [7:0]  io_weight_win_33_512,
  input  [7:0]  io_weight_win_33_513,
  input  [7:0]  io_weight_win_33_514,
  input  [7:0]  io_weight_win_33_515,
  input  [7:0]  io_weight_win_33_516,
  input  [7:0]  io_weight_win_33_517,
  input  [7:0]  io_weight_win_33_518,
  input  [7:0]  io_weight_win_33_519,
  input  [7:0]  io_weight_win_33_520,
  input  [7:0]  io_weight_win_33_521,
  input  [7:0]  io_weight_win_33_522,
  input  [7:0]  io_weight_win_33_523,
  input  [7:0]  io_weight_win_33_524,
  input  [7:0]  io_weight_win_33_525,
  input  [7:0]  io_weight_win_33_526,
  input  [7:0]  io_weight_win_33_527,
  input  [7:0]  io_weight_win_33_528,
  input  [7:0]  io_weight_win_33_529,
  input  [7:0]  io_weight_win_33_530,
  input  [7:0]  io_weight_win_33_531,
  input  [7:0]  io_weight_win_33_532,
  input  [7:0]  io_weight_win_33_533,
  input  [7:0]  io_weight_win_33_534,
  input  [7:0]  io_weight_win_33_535,
  input  [7:0]  io_weight_win_33_536,
  input  [7:0]  io_weight_win_33_537,
  input  [7:0]  io_weight_win_33_538,
  input  [7:0]  io_weight_win_33_539,
  input  [7:0]  io_weight_win_33_540,
  input  [7:0]  io_weight_win_33_541,
  input  [7:0]  io_weight_win_33_542,
  input  [7:0]  io_weight_win_33_543,
  input  [7:0]  io_weight_win_33_544,
  input  [7:0]  io_weight_win_33_545,
  input  [7:0]  io_weight_win_33_546,
  input  [7:0]  io_weight_win_33_547,
  input  [7:0]  io_weight_win_33_548,
  input  [7:0]  io_weight_win_33_549,
  input  [7:0]  io_weight_win_33_550,
  input  [7:0]  io_weight_win_33_551,
  input  [7:0]  io_weight_win_33_552,
  input  [7:0]  io_weight_win_33_553,
  input  [7:0]  io_weight_win_33_554,
  input  [7:0]  io_weight_win_33_555,
  input  [7:0]  io_weight_win_33_556,
  input  [7:0]  io_weight_win_33_557,
  input  [7:0]  io_weight_win_33_558,
  input  [7:0]  io_weight_win_33_559,
  input  [7:0]  io_weight_win_33_560,
  input  [7:0]  io_weight_win_33_561,
  input  [7:0]  io_weight_win_33_562,
  input  [7:0]  io_weight_win_33_563,
  input  [7:0]  io_weight_win_33_564,
  input  [7:0]  io_weight_win_33_565,
  input  [7:0]  io_weight_win_33_566,
  input  [7:0]  io_weight_win_33_567,
  input  [7:0]  io_weight_win_33_568,
  input  [7:0]  io_weight_win_33_569,
  input  [7:0]  io_weight_win_33_570,
  input  [7:0]  io_weight_win_33_571,
  input  [7:0]  io_weight_win_33_572,
  input  [7:0]  io_weight_win_33_573,
  input  [7:0]  io_weight_win_33_574,
  input  [7:0]  io_weight_win_33_575,
  input  [17:0] io_bias_data_0,
  input  [17:0] io_bias_data_1,
  input  [17:0] io_bias_data_2,
  input  [17:0] io_bias_data_3,
  input  [17:0] io_bias_data_4,
  input  [17:0] io_bias_data_5,
  input  [17:0] io_bias_data_6,
  input  [17:0] io_bias_data_7,
  input         io_bias_valid,
  output [17:0] io_conv_o_0,
  output [17:0] io_conv_o_1,
  output [17:0] io_conv_o_2,
  output [17:0] io_conv_o_3,
  output [17:0] io_conv_o_4,
  output [17:0] io_conv_o_5,
  output [17:0] io_conv_o_6,
  output [17:0] io_conv_o_7
);
  wire  conv_unit_0_clock; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_ifm_win_33_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch1_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_0_io_weight_win_33_ch2_71; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_0_io_bias1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_0_io_bias2; // @[Conv.scala 18:47]
  wire  conv_unit_0_io_bias_valid; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_0_io_o_conv_ch1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_0_io_o_conv_ch2; // @[Conv.scala 18:47]
  wire  conv_unit_1_clock; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_ifm_win_33_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch1_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_1_io_weight_win_33_ch2_71; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_1_io_bias1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_1_io_bias2; // @[Conv.scala 18:47]
  wire  conv_unit_1_io_bias_valid; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_1_io_o_conv_ch1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_1_io_o_conv_ch2; // @[Conv.scala 18:47]
  wire  conv_unit_2_clock; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_ifm_win_33_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch1_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_2_io_weight_win_33_ch2_71; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_2_io_bias1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_2_io_bias2; // @[Conv.scala 18:47]
  wire  conv_unit_2_io_bias_valid; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_2_io_o_conv_ch1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_2_io_o_conv_ch2; // @[Conv.scala 18:47]
  wire  conv_unit_3_clock; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_ifm_win_33_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch1_71; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_0; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_1; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_2; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_3; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_4; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_5; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_6; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_7; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_8; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_9; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_10; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_11; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_12; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_13; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_14; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_15; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_16; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_17; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_18; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_19; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_20; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_21; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_22; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_23; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_24; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_25; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_26; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_27; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_28; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_29; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_30; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_31; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_32; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_33; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_34; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_35; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_36; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_37; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_38; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_39; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_40; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_41; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_42; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_43; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_44; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_45; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_46; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_47; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_48; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_49; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_50; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_51; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_52; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_53; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_54; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_55; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_56; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_57; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_58; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_59; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_60; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_61; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_62; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_63; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_64; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_65; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_66; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_67; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_68; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_69; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_70; // @[Conv.scala 18:47]
  wire [7:0] conv_unit_3_io_weight_win_33_ch2_71; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_3_io_bias1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_3_io_bias2; // @[Conv.scala 18:47]
  wire  conv_unit_3_io_bias_valid; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_3_io_o_conv_ch1; // @[Conv.scala 18:47]
  wire [17:0] conv_unit_3_io_o_conv_ch2; // @[Conv.scala 18:47]
  conv_unit conv_unit_0 ( // @[Conv.scala 18:47]
    .clock(conv_unit_0_clock),
    .io_ifm_win_33_0(conv_unit_0_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_unit_0_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_unit_0_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_unit_0_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_unit_0_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_unit_0_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_unit_0_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_unit_0_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_unit_0_io_ifm_win_33_8),
    .io_ifm_win_33_9(conv_unit_0_io_ifm_win_33_9),
    .io_ifm_win_33_10(conv_unit_0_io_ifm_win_33_10),
    .io_ifm_win_33_11(conv_unit_0_io_ifm_win_33_11),
    .io_ifm_win_33_12(conv_unit_0_io_ifm_win_33_12),
    .io_ifm_win_33_13(conv_unit_0_io_ifm_win_33_13),
    .io_ifm_win_33_14(conv_unit_0_io_ifm_win_33_14),
    .io_ifm_win_33_15(conv_unit_0_io_ifm_win_33_15),
    .io_ifm_win_33_16(conv_unit_0_io_ifm_win_33_16),
    .io_ifm_win_33_17(conv_unit_0_io_ifm_win_33_17),
    .io_ifm_win_33_18(conv_unit_0_io_ifm_win_33_18),
    .io_ifm_win_33_19(conv_unit_0_io_ifm_win_33_19),
    .io_ifm_win_33_20(conv_unit_0_io_ifm_win_33_20),
    .io_ifm_win_33_21(conv_unit_0_io_ifm_win_33_21),
    .io_ifm_win_33_22(conv_unit_0_io_ifm_win_33_22),
    .io_ifm_win_33_23(conv_unit_0_io_ifm_win_33_23),
    .io_ifm_win_33_24(conv_unit_0_io_ifm_win_33_24),
    .io_ifm_win_33_25(conv_unit_0_io_ifm_win_33_25),
    .io_ifm_win_33_26(conv_unit_0_io_ifm_win_33_26),
    .io_ifm_win_33_27(conv_unit_0_io_ifm_win_33_27),
    .io_ifm_win_33_28(conv_unit_0_io_ifm_win_33_28),
    .io_ifm_win_33_29(conv_unit_0_io_ifm_win_33_29),
    .io_ifm_win_33_30(conv_unit_0_io_ifm_win_33_30),
    .io_ifm_win_33_31(conv_unit_0_io_ifm_win_33_31),
    .io_ifm_win_33_32(conv_unit_0_io_ifm_win_33_32),
    .io_ifm_win_33_33(conv_unit_0_io_ifm_win_33_33),
    .io_ifm_win_33_34(conv_unit_0_io_ifm_win_33_34),
    .io_ifm_win_33_35(conv_unit_0_io_ifm_win_33_35),
    .io_ifm_win_33_36(conv_unit_0_io_ifm_win_33_36),
    .io_ifm_win_33_37(conv_unit_0_io_ifm_win_33_37),
    .io_ifm_win_33_38(conv_unit_0_io_ifm_win_33_38),
    .io_ifm_win_33_39(conv_unit_0_io_ifm_win_33_39),
    .io_ifm_win_33_40(conv_unit_0_io_ifm_win_33_40),
    .io_ifm_win_33_41(conv_unit_0_io_ifm_win_33_41),
    .io_ifm_win_33_42(conv_unit_0_io_ifm_win_33_42),
    .io_ifm_win_33_43(conv_unit_0_io_ifm_win_33_43),
    .io_ifm_win_33_44(conv_unit_0_io_ifm_win_33_44),
    .io_ifm_win_33_45(conv_unit_0_io_ifm_win_33_45),
    .io_ifm_win_33_46(conv_unit_0_io_ifm_win_33_46),
    .io_ifm_win_33_47(conv_unit_0_io_ifm_win_33_47),
    .io_ifm_win_33_48(conv_unit_0_io_ifm_win_33_48),
    .io_ifm_win_33_49(conv_unit_0_io_ifm_win_33_49),
    .io_ifm_win_33_50(conv_unit_0_io_ifm_win_33_50),
    .io_ifm_win_33_51(conv_unit_0_io_ifm_win_33_51),
    .io_ifm_win_33_52(conv_unit_0_io_ifm_win_33_52),
    .io_ifm_win_33_53(conv_unit_0_io_ifm_win_33_53),
    .io_ifm_win_33_54(conv_unit_0_io_ifm_win_33_54),
    .io_ifm_win_33_55(conv_unit_0_io_ifm_win_33_55),
    .io_ifm_win_33_56(conv_unit_0_io_ifm_win_33_56),
    .io_ifm_win_33_57(conv_unit_0_io_ifm_win_33_57),
    .io_ifm_win_33_58(conv_unit_0_io_ifm_win_33_58),
    .io_ifm_win_33_59(conv_unit_0_io_ifm_win_33_59),
    .io_ifm_win_33_60(conv_unit_0_io_ifm_win_33_60),
    .io_ifm_win_33_61(conv_unit_0_io_ifm_win_33_61),
    .io_ifm_win_33_62(conv_unit_0_io_ifm_win_33_62),
    .io_ifm_win_33_63(conv_unit_0_io_ifm_win_33_63),
    .io_ifm_win_33_64(conv_unit_0_io_ifm_win_33_64),
    .io_ifm_win_33_65(conv_unit_0_io_ifm_win_33_65),
    .io_ifm_win_33_66(conv_unit_0_io_ifm_win_33_66),
    .io_ifm_win_33_67(conv_unit_0_io_ifm_win_33_67),
    .io_ifm_win_33_68(conv_unit_0_io_ifm_win_33_68),
    .io_ifm_win_33_69(conv_unit_0_io_ifm_win_33_69),
    .io_ifm_win_33_70(conv_unit_0_io_ifm_win_33_70),
    .io_ifm_win_33_71(conv_unit_0_io_ifm_win_33_71),
    .io_weight_win_33_ch1_0(conv_unit_0_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_unit_0_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_unit_0_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_unit_0_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_unit_0_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_unit_0_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_unit_0_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_unit_0_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_unit_0_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch1_9(conv_unit_0_io_weight_win_33_ch1_9),
    .io_weight_win_33_ch1_10(conv_unit_0_io_weight_win_33_ch1_10),
    .io_weight_win_33_ch1_11(conv_unit_0_io_weight_win_33_ch1_11),
    .io_weight_win_33_ch1_12(conv_unit_0_io_weight_win_33_ch1_12),
    .io_weight_win_33_ch1_13(conv_unit_0_io_weight_win_33_ch1_13),
    .io_weight_win_33_ch1_14(conv_unit_0_io_weight_win_33_ch1_14),
    .io_weight_win_33_ch1_15(conv_unit_0_io_weight_win_33_ch1_15),
    .io_weight_win_33_ch1_16(conv_unit_0_io_weight_win_33_ch1_16),
    .io_weight_win_33_ch1_17(conv_unit_0_io_weight_win_33_ch1_17),
    .io_weight_win_33_ch1_18(conv_unit_0_io_weight_win_33_ch1_18),
    .io_weight_win_33_ch1_19(conv_unit_0_io_weight_win_33_ch1_19),
    .io_weight_win_33_ch1_20(conv_unit_0_io_weight_win_33_ch1_20),
    .io_weight_win_33_ch1_21(conv_unit_0_io_weight_win_33_ch1_21),
    .io_weight_win_33_ch1_22(conv_unit_0_io_weight_win_33_ch1_22),
    .io_weight_win_33_ch1_23(conv_unit_0_io_weight_win_33_ch1_23),
    .io_weight_win_33_ch1_24(conv_unit_0_io_weight_win_33_ch1_24),
    .io_weight_win_33_ch1_25(conv_unit_0_io_weight_win_33_ch1_25),
    .io_weight_win_33_ch1_26(conv_unit_0_io_weight_win_33_ch1_26),
    .io_weight_win_33_ch1_27(conv_unit_0_io_weight_win_33_ch1_27),
    .io_weight_win_33_ch1_28(conv_unit_0_io_weight_win_33_ch1_28),
    .io_weight_win_33_ch1_29(conv_unit_0_io_weight_win_33_ch1_29),
    .io_weight_win_33_ch1_30(conv_unit_0_io_weight_win_33_ch1_30),
    .io_weight_win_33_ch1_31(conv_unit_0_io_weight_win_33_ch1_31),
    .io_weight_win_33_ch1_32(conv_unit_0_io_weight_win_33_ch1_32),
    .io_weight_win_33_ch1_33(conv_unit_0_io_weight_win_33_ch1_33),
    .io_weight_win_33_ch1_34(conv_unit_0_io_weight_win_33_ch1_34),
    .io_weight_win_33_ch1_35(conv_unit_0_io_weight_win_33_ch1_35),
    .io_weight_win_33_ch1_36(conv_unit_0_io_weight_win_33_ch1_36),
    .io_weight_win_33_ch1_37(conv_unit_0_io_weight_win_33_ch1_37),
    .io_weight_win_33_ch1_38(conv_unit_0_io_weight_win_33_ch1_38),
    .io_weight_win_33_ch1_39(conv_unit_0_io_weight_win_33_ch1_39),
    .io_weight_win_33_ch1_40(conv_unit_0_io_weight_win_33_ch1_40),
    .io_weight_win_33_ch1_41(conv_unit_0_io_weight_win_33_ch1_41),
    .io_weight_win_33_ch1_42(conv_unit_0_io_weight_win_33_ch1_42),
    .io_weight_win_33_ch1_43(conv_unit_0_io_weight_win_33_ch1_43),
    .io_weight_win_33_ch1_44(conv_unit_0_io_weight_win_33_ch1_44),
    .io_weight_win_33_ch1_45(conv_unit_0_io_weight_win_33_ch1_45),
    .io_weight_win_33_ch1_46(conv_unit_0_io_weight_win_33_ch1_46),
    .io_weight_win_33_ch1_47(conv_unit_0_io_weight_win_33_ch1_47),
    .io_weight_win_33_ch1_48(conv_unit_0_io_weight_win_33_ch1_48),
    .io_weight_win_33_ch1_49(conv_unit_0_io_weight_win_33_ch1_49),
    .io_weight_win_33_ch1_50(conv_unit_0_io_weight_win_33_ch1_50),
    .io_weight_win_33_ch1_51(conv_unit_0_io_weight_win_33_ch1_51),
    .io_weight_win_33_ch1_52(conv_unit_0_io_weight_win_33_ch1_52),
    .io_weight_win_33_ch1_53(conv_unit_0_io_weight_win_33_ch1_53),
    .io_weight_win_33_ch1_54(conv_unit_0_io_weight_win_33_ch1_54),
    .io_weight_win_33_ch1_55(conv_unit_0_io_weight_win_33_ch1_55),
    .io_weight_win_33_ch1_56(conv_unit_0_io_weight_win_33_ch1_56),
    .io_weight_win_33_ch1_57(conv_unit_0_io_weight_win_33_ch1_57),
    .io_weight_win_33_ch1_58(conv_unit_0_io_weight_win_33_ch1_58),
    .io_weight_win_33_ch1_59(conv_unit_0_io_weight_win_33_ch1_59),
    .io_weight_win_33_ch1_60(conv_unit_0_io_weight_win_33_ch1_60),
    .io_weight_win_33_ch1_61(conv_unit_0_io_weight_win_33_ch1_61),
    .io_weight_win_33_ch1_62(conv_unit_0_io_weight_win_33_ch1_62),
    .io_weight_win_33_ch1_63(conv_unit_0_io_weight_win_33_ch1_63),
    .io_weight_win_33_ch1_64(conv_unit_0_io_weight_win_33_ch1_64),
    .io_weight_win_33_ch1_65(conv_unit_0_io_weight_win_33_ch1_65),
    .io_weight_win_33_ch1_66(conv_unit_0_io_weight_win_33_ch1_66),
    .io_weight_win_33_ch1_67(conv_unit_0_io_weight_win_33_ch1_67),
    .io_weight_win_33_ch1_68(conv_unit_0_io_weight_win_33_ch1_68),
    .io_weight_win_33_ch1_69(conv_unit_0_io_weight_win_33_ch1_69),
    .io_weight_win_33_ch1_70(conv_unit_0_io_weight_win_33_ch1_70),
    .io_weight_win_33_ch1_71(conv_unit_0_io_weight_win_33_ch1_71),
    .io_weight_win_33_ch2_0(conv_unit_0_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_unit_0_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_unit_0_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_unit_0_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_unit_0_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_unit_0_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_unit_0_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_unit_0_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_unit_0_io_weight_win_33_ch2_8),
    .io_weight_win_33_ch2_9(conv_unit_0_io_weight_win_33_ch2_9),
    .io_weight_win_33_ch2_10(conv_unit_0_io_weight_win_33_ch2_10),
    .io_weight_win_33_ch2_11(conv_unit_0_io_weight_win_33_ch2_11),
    .io_weight_win_33_ch2_12(conv_unit_0_io_weight_win_33_ch2_12),
    .io_weight_win_33_ch2_13(conv_unit_0_io_weight_win_33_ch2_13),
    .io_weight_win_33_ch2_14(conv_unit_0_io_weight_win_33_ch2_14),
    .io_weight_win_33_ch2_15(conv_unit_0_io_weight_win_33_ch2_15),
    .io_weight_win_33_ch2_16(conv_unit_0_io_weight_win_33_ch2_16),
    .io_weight_win_33_ch2_17(conv_unit_0_io_weight_win_33_ch2_17),
    .io_weight_win_33_ch2_18(conv_unit_0_io_weight_win_33_ch2_18),
    .io_weight_win_33_ch2_19(conv_unit_0_io_weight_win_33_ch2_19),
    .io_weight_win_33_ch2_20(conv_unit_0_io_weight_win_33_ch2_20),
    .io_weight_win_33_ch2_21(conv_unit_0_io_weight_win_33_ch2_21),
    .io_weight_win_33_ch2_22(conv_unit_0_io_weight_win_33_ch2_22),
    .io_weight_win_33_ch2_23(conv_unit_0_io_weight_win_33_ch2_23),
    .io_weight_win_33_ch2_24(conv_unit_0_io_weight_win_33_ch2_24),
    .io_weight_win_33_ch2_25(conv_unit_0_io_weight_win_33_ch2_25),
    .io_weight_win_33_ch2_26(conv_unit_0_io_weight_win_33_ch2_26),
    .io_weight_win_33_ch2_27(conv_unit_0_io_weight_win_33_ch2_27),
    .io_weight_win_33_ch2_28(conv_unit_0_io_weight_win_33_ch2_28),
    .io_weight_win_33_ch2_29(conv_unit_0_io_weight_win_33_ch2_29),
    .io_weight_win_33_ch2_30(conv_unit_0_io_weight_win_33_ch2_30),
    .io_weight_win_33_ch2_31(conv_unit_0_io_weight_win_33_ch2_31),
    .io_weight_win_33_ch2_32(conv_unit_0_io_weight_win_33_ch2_32),
    .io_weight_win_33_ch2_33(conv_unit_0_io_weight_win_33_ch2_33),
    .io_weight_win_33_ch2_34(conv_unit_0_io_weight_win_33_ch2_34),
    .io_weight_win_33_ch2_35(conv_unit_0_io_weight_win_33_ch2_35),
    .io_weight_win_33_ch2_36(conv_unit_0_io_weight_win_33_ch2_36),
    .io_weight_win_33_ch2_37(conv_unit_0_io_weight_win_33_ch2_37),
    .io_weight_win_33_ch2_38(conv_unit_0_io_weight_win_33_ch2_38),
    .io_weight_win_33_ch2_39(conv_unit_0_io_weight_win_33_ch2_39),
    .io_weight_win_33_ch2_40(conv_unit_0_io_weight_win_33_ch2_40),
    .io_weight_win_33_ch2_41(conv_unit_0_io_weight_win_33_ch2_41),
    .io_weight_win_33_ch2_42(conv_unit_0_io_weight_win_33_ch2_42),
    .io_weight_win_33_ch2_43(conv_unit_0_io_weight_win_33_ch2_43),
    .io_weight_win_33_ch2_44(conv_unit_0_io_weight_win_33_ch2_44),
    .io_weight_win_33_ch2_45(conv_unit_0_io_weight_win_33_ch2_45),
    .io_weight_win_33_ch2_46(conv_unit_0_io_weight_win_33_ch2_46),
    .io_weight_win_33_ch2_47(conv_unit_0_io_weight_win_33_ch2_47),
    .io_weight_win_33_ch2_48(conv_unit_0_io_weight_win_33_ch2_48),
    .io_weight_win_33_ch2_49(conv_unit_0_io_weight_win_33_ch2_49),
    .io_weight_win_33_ch2_50(conv_unit_0_io_weight_win_33_ch2_50),
    .io_weight_win_33_ch2_51(conv_unit_0_io_weight_win_33_ch2_51),
    .io_weight_win_33_ch2_52(conv_unit_0_io_weight_win_33_ch2_52),
    .io_weight_win_33_ch2_53(conv_unit_0_io_weight_win_33_ch2_53),
    .io_weight_win_33_ch2_54(conv_unit_0_io_weight_win_33_ch2_54),
    .io_weight_win_33_ch2_55(conv_unit_0_io_weight_win_33_ch2_55),
    .io_weight_win_33_ch2_56(conv_unit_0_io_weight_win_33_ch2_56),
    .io_weight_win_33_ch2_57(conv_unit_0_io_weight_win_33_ch2_57),
    .io_weight_win_33_ch2_58(conv_unit_0_io_weight_win_33_ch2_58),
    .io_weight_win_33_ch2_59(conv_unit_0_io_weight_win_33_ch2_59),
    .io_weight_win_33_ch2_60(conv_unit_0_io_weight_win_33_ch2_60),
    .io_weight_win_33_ch2_61(conv_unit_0_io_weight_win_33_ch2_61),
    .io_weight_win_33_ch2_62(conv_unit_0_io_weight_win_33_ch2_62),
    .io_weight_win_33_ch2_63(conv_unit_0_io_weight_win_33_ch2_63),
    .io_weight_win_33_ch2_64(conv_unit_0_io_weight_win_33_ch2_64),
    .io_weight_win_33_ch2_65(conv_unit_0_io_weight_win_33_ch2_65),
    .io_weight_win_33_ch2_66(conv_unit_0_io_weight_win_33_ch2_66),
    .io_weight_win_33_ch2_67(conv_unit_0_io_weight_win_33_ch2_67),
    .io_weight_win_33_ch2_68(conv_unit_0_io_weight_win_33_ch2_68),
    .io_weight_win_33_ch2_69(conv_unit_0_io_weight_win_33_ch2_69),
    .io_weight_win_33_ch2_70(conv_unit_0_io_weight_win_33_ch2_70),
    .io_weight_win_33_ch2_71(conv_unit_0_io_weight_win_33_ch2_71),
    .io_bias1(conv_unit_0_io_bias1),
    .io_bias2(conv_unit_0_io_bias2),
    .io_bias_valid(conv_unit_0_io_bias_valid),
    .io_o_conv_ch1(conv_unit_0_io_o_conv_ch1),
    .io_o_conv_ch2(conv_unit_0_io_o_conv_ch2)
  );
  conv_unit conv_unit_1 ( // @[Conv.scala 18:47]
    .clock(conv_unit_1_clock),
    .io_ifm_win_33_0(conv_unit_1_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_unit_1_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_unit_1_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_unit_1_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_unit_1_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_unit_1_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_unit_1_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_unit_1_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_unit_1_io_ifm_win_33_8),
    .io_ifm_win_33_9(conv_unit_1_io_ifm_win_33_9),
    .io_ifm_win_33_10(conv_unit_1_io_ifm_win_33_10),
    .io_ifm_win_33_11(conv_unit_1_io_ifm_win_33_11),
    .io_ifm_win_33_12(conv_unit_1_io_ifm_win_33_12),
    .io_ifm_win_33_13(conv_unit_1_io_ifm_win_33_13),
    .io_ifm_win_33_14(conv_unit_1_io_ifm_win_33_14),
    .io_ifm_win_33_15(conv_unit_1_io_ifm_win_33_15),
    .io_ifm_win_33_16(conv_unit_1_io_ifm_win_33_16),
    .io_ifm_win_33_17(conv_unit_1_io_ifm_win_33_17),
    .io_ifm_win_33_18(conv_unit_1_io_ifm_win_33_18),
    .io_ifm_win_33_19(conv_unit_1_io_ifm_win_33_19),
    .io_ifm_win_33_20(conv_unit_1_io_ifm_win_33_20),
    .io_ifm_win_33_21(conv_unit_1_io_ifm_win_33_21),
    .io_ifm_win_33_22(conv_unit_1_io_ifm_win_33_22),
    .io_ifm_win_33_23(conv_unit_1_io_ifm_win_33_23),
    .io_ifm_win_33_24(conv_unit_1_io_ifm_win_33_24),
    .io_ifm_win_33_25(conv_unit_1_io_ifm_win_33_25),
    .io_ifm_win_33_26(conv_unit_1_io_ifm_win_33_26),
    .io_ifm_win_33_27(conv_unit_1_io_ifm_win_33_27),
    .io_ifm_win_33_28(conv_unit_1_io_ifm_win_33_28),
    .io_ifm_win_33_29(conv_unit_1_io_ifm_win_33_29),
    .io_ifm_win_33_30(conv_unit_1_io_ifm_win_33_30),
    .io_ifm_win_33_31(conv_unit_1_io_ifm_win_33_31),
    .io_ifm_win_33_32(conv_unit_1_io_ifm_win_33_32),
    .io_ifm_win_33_33(conv_unit_1_io_ifm_win_33_33),
    .io_ifm_win_33_34(conv_unit_1_io_ifm_win_33_34),
    .io_ifm_win_33_35(conv_unit_1_io_ifm_win_33_35),
    .io_ifm_win_33_36(conv_unit_1_io_ifm_win_33_36),
    .io_ifm_win_33_37(conv_unit_1_io_ifm_win_33_37),
    .io_ifm_win_33_38(conv_unit_1_io_ifm_win_33_38),
    .io_ifm_win_33_39(conv_unit_1_io_ifm_win_33_39),
    .io_ifm_win_33_40(conv_unit_1_io_ifm_win_33_40),
    .io_ifm_win_33_41(conv_unit_1_io_ifm_win_33_41),
    .io_ifm_win_33_42(conv_unit_1_io_ifm_win_33_42),
    .io_ifm_win_33_43(conv_unit_1_io_ifm_win_33_43),
    .io_ifm_win_33_44(conv_unit_1_io_ifm_win_33_44),
    .io_ifm_win_33_45(conv_unit_1_io_ifm_win_33_45),
    .io_ifm_win_33_46(conv_unit_1_io_ifm_win_33_46),
    .io_ifm_win_33_47(conv_unit_1_io_ifm_win_33_47),
    .io_ifm_win_33_48(conv_unit_1_io_ifm_win_33_48),
    .io_ifm_win_33_49(conv_unit_1_io_ifm_win_33_49),
    .io_ifm_win_33_50(conv_unit_1_io_ifm_win_33_50),
    .io_ifm_win_33_51(conv_unit_1_io_ifm_win_33_51),
    .io_ifm_win_33_52(conv_unit_1_io_ifm_win_33_52),
    .io_ifm_win_33_53(conv_unit_1_io_ifm_win_33_53),
    .io_ifm_win_33_54(conv_unit_1_io_ifm_win_33_54),
    .io_ifm_win_33_55(conv_unit_1_io_ifm_win_33_55),
    .io_ifm_win_33_56(conv_unit_1_io_ifm_win_33_56),
    .io_ifm_win_33_57(conv_unit_1_io_ifm_win_33_57),
    .io_ifm_win_33_58(conv_unit_1_io_ifm_win_33_58),
    .io_ifm_win_33_59(conv_unit_1_io_ifm_win_33_59),
    .io_ifm_win_33_60(conv_unit_1_io_ifm_win_33_60),
    .io_ifm_win_33_61(conv_unit_1_io_ifm_win_33_61),
    .io_ifm_win_33_62(conv_unit_1_io_ifm_win_33_62),
    .io_ifm_win_33_63(conv_unit_1_io_ifm_win_33_63),
    .io_ifm_win_33_64(conv_unit_1_io_ifm_win_33_64),
    .io_ifm_win_33_65(conv_unit_1_io_ifm_win_33_65),
    .io_ifm_win_33_66(conv_unit_1_io_ifm_win_33_66),
    .io_ifm_win_33_67(conv_unit_1_io_ifm_win_33_67),
    .io_ifm_win_33_68(conv_unit_1_io_ifm_win_33_68),
    .io_ifm_win_33_69(conv_unit_1_io_ifm_win_33_69),
    .io_ifm_win_33_70(conv_unit_1_io_ifm_win_33_70),
    .io_ifm_win_33_71(conv_unit_1_io_ifm_win_33_71),
    .io_weight_win_33_ch1_0(conv_unit_1_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_unit_1_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_unit_1_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_unit_1_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_unit_1_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_unit_1_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_unit_1_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_unit_1_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_unit_1_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch1_9(conv_unit_1_io_weight_win_33_ch1_9),
    .io_weight_win_33_ch1_10(conv_unit_1_io_weight_win_33_ch1_10),
    .io_weight_win_33_ch1_11(conv_unit_1_io_weight_win_33_ch1_11),
    .io_weight_win_33_ch1_12(conv_unit_1_io_weight_win_33_ch1_12),
    .io_weight_win_33_ch1_13(conv_unit_1_io_weight_win_33_ch1_13),
    .io_weight_win_33_ch1_14(conv_unit_1_io_weight_win_33_ch1_14),
    .io_weight_win_33_ch1_15(conv_unit_1_io_weight_win_33_ch1_15),
    .io_weight_win_33_ch1_16(conv_unit_1_io_weight_win_33_ch1_16),
    .io_weight_win_33_ch1_17(conv_unit_1_io_weight_win_33_ch1_17),
    .io_weight_win_33_ch1_18(conv_unit_1_io_weight_win_33_ch1_18),
    .io_weight_win_33_ch1_19(conv_unit_1_io_weight_win_33_ch1_19),
    .io_weight_win_33_ch1_20(conv_unit_1_io_weight_win_33_ch1_20),
    .io_weight_win_33_ch1_21(conv_unit_1_io_weight_win_33_ch1_21),
    .io_weight_win_33_ch1_22(conv_unit_1_io_weight_win_33_ch1_22),
    .io_weight_win_33_ch1_23(conv_unit_1_io_weight_win_33_ch1_23),
    .io_weight_win_33_ch1_24(conv_unit_1_io_weight_win_33_ch1_24),
    .io_weight_win_33_ch1_25(conv_unit_1_io_weight_win_33_ch1_25),
    .io_weight_win_33_ch1_26(conv_unit_1_io_weight_win_33_ch1_26),
    .io_weight_win_33_ch1_27(conv_unit_1_io_weight_win_33_ch1_27),
    .io_weight_win_33_ch1_28(conv_unit_1_io_weight_win_33_ch1_28),
    .io_weight_win_33_ch1_29(conv_unit_1_io_weight_win_33_ch1_29),
    .io_weight_win_33_ch1_30(conv_unit_1_io_weight_win_33_ch1_30),
    .io_weight_win_33_ch1_31(conv_unit_1_io_weight_win_33_ch1_31),
    .io_weight_win_33_ch1_32(conv_unit_1_io_weight_win_33_ch1_32),
    .io_weight_win_33_ch1_33(conv_unit_1_io_weight_win_33_ch1_33),
    .io_weight_win_33_ch1_34(conv_unit_1_io_weight_win_33_ch1_34),
    .io_weight_win_33_ch1_35(conv_unit_1_io_weight_win_33_ch1_35),
    .io_weight_win_33_ch1_36(conv_unit_1_io_weight_win_33_ch1_36),
    .io_weight_win_33_ch1_37(conv_unit_1_io_weight_win_33_ch1_37),
    .io_weight_win_33_ch1_38(conv_unit_1_io_weight_win_33_ch1_38),
    .io_weight_win_33_ch1_39(conv_unit_1_io_weight_win_33_ch1_39),
    .io_weight_win_33_ch1_40(conv_unit_1_io_weight_win_33_ch1_40),
    .io_weight_win_33_ch1_41(conv_unit_1_io_weight_win_33_ch1_41),
    .io_weight_win_33_ch1_42(conv_unit_1_io_weight_win_33_ch1_42),
    .io_weight_win_33_ch1_43(conv_unit_1_io_weight_win_33_ch1_43),
    .io_weight_win_33_ch1_44(conv_unit_1_io_weight_win_33_ch1_44),
    .io_weight_win_33_ch1_45(conv_unit_1_io_weight_win_33_ch1_45),
    .io_weight_win_33_ch1_46(conv_unit_1_io_weight_win_33_ch1_46),
    .io_weight_win_33_ch1_47(conv_unit_1_io_weight_win_33_ch1_47),
    .io_weight_win_33_ch1_48(conv_unit_1_io_weight_win_33_ch1_48),
    .io_weight_win_33_ch1_49(conv_unit_1_io_weight_win_33_ch1_49),
    .io_weight_win_33_ch1_50(conv_unit_1_io_weight_win_33_ch1_50),
    .io_weight_win_33_ch1_51(conv_unit_1_io_weight_win_33_ch1_51),
    .io_weight_win_33_ch1_52(conv_unit_1_io_weight_win_33_ch1_52),
    .io_weight_win_33_ch1_53(conv_unit_1_io_weight_win_33_ch1_53),
    .io_weight_win_33_ch1_54(conv_unit_1_io_weight_win_33_ch1_54),
    .io_weight_win_33_ch1_55(conv_unit_1_io_weight_win_33_ch1_55),
    .io_weight_win_33_ch1_56(conv_unit_1_io_weight_win_33_ch1_56),
    .io_weight_win_33_ch1_57(conv_unit_1_io_weight_win_33_ch1_57),
    .io_weight_win_33_ch1_58(conv_unit_1_io_weight_win_33_ch1_58),
    .io_weight_win_33_ch1_59(conv_unit_1_io_weight_win_33_ch1_59),
    .io_weight_win_33_ch1_60(conv_unit_1_io_weight_win_33_ch1_60),
    .io_weight_win_33_ch1_61(conv_unit_1_io_weight_win_33_ch1_61),
    .io_weight_win_33_ch1_62(conv_unit_1_io_weight_win_33_ch1_62),
    .io_weight_win_33_ch1_63(conv_unit_1_io_weight_win_33_ch1_63),
    .io_weight_win_33_ch1_64(conv_unit_1_io_weight_win_33_ch1_64),
    .io_weight_win_33_ch1_65(conv_unit_1_io_weight_win_33_ch1_65),
    .io_weight_win_33_ch1_66(conv_unit_1_io_weight_win_33_ch1_66),
    .io_weight_win_33_ch1_67(conv_unit_1_io_weight_win_33_ch1_67),
    .io_weight_win_33_ch1_68(conv_unit_1_io_weight_win_33_ch1_68),
    .io_weight_win_33_ch1_69(conv_unit_1_io_weight_win_33_ch1_69),
    .io_weight_win_33_ch1_70(conv_unit_1_io_weight_win_33_ch1_70),
    .io_weight_win_33_ch1_71(conv_unit_1_io_weight_win_33_ch1_71),
    .io_weight_win_33_ch2_0(conv_unit_1_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_unit_1_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_unit_1_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_unit_1_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_unit_1_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_unit_1_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_unit_1_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_unit_1_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_unit_1_io_weight_win_33_ch2_8),
    .io_weight_win_33_ch2_9(conv_unit_1_io_weight_win_33_ch2_9),
    .io_weight_win_33_ch2_10(conv_unit_1_io_weight_win_33_ch2_10),
    .io_weight_win_33_ch2_11(conv_unit_1_io_weight_win_33_ch2_11),
    .io_weight_win_33_ch2_12(conv_unit_1_io_weight_win_33_ch2_12),
    .io_weight_win_33_ch2_13(conv_unit_1_io_weight_win_33_ch2_13),
    .io_weight_win_33_ch2_14(conv_unit_1_io_weight_win_33_ch2_14),
    .io_weight_win_33_ch2_15(conv_unit_1_io_weight_win_33_ch2_15),
    .io_weight_win_33_ch2_16(conv_unit_1_io_weight_win_33_ch2_16),
    .io_weight_win_33_ch2_17(conv_unit_1_io_weight_win_33_ch2_17),
    .io_weight_win_33_ch2_18(conv_unit_1_io_weight_win_33_ch2_18),
    .io_weight_win_33_ch2_19(conv_unit_1_io_weight_win_33_ch2_19),
    .io_weight_win_33_ch2_20(conv_unit_1_io_weight_win_33_ch2_20),
    .io_weight_win_33_ch2_21(conv_unit_1_io_weight_win_33_ch2_21),
    .io_weight_win_33_ch2_22(conv_unit_1_io_weight_win_33_ch2_22),
    .io_weight_win_33_ch2_23(conv_unit_1_io_weight_win_33_ch2_23),
    .io_weight_win_33_ch2_24(conv_unit_1_io_weight_win_33_ch2_24),
    .io_weight_win_33_ch2_25(conv_unit_1_io_weight_win_33_ch2_25),
    .io_weight_win_33_ch2_26(conv_unit_1_io_weight_win_33_ch2_26),
    .io_weight_win_33_ch2_27(conv_unit_1_io_weight_win_33_ch2_27),
    .io_weight_win_33_ch2_28(conv_unit_1_io_weight_win_33_ch2_28),
    .io_weight_win_33_ch2_29(conv_unit_1_io_weight_win_33_ch2_29),
    .io_weight_win_33_ch2_30(conv_unit_1_io_weight_win_33_ch2_30),
    .io_weight_win_33_ch2_31(conv_unit_1_io_weight_win_33_ch2_31),
    .io_weight_win_33_ch2_32(conv_unit_1_io_weight_win_33_ch2_32),
    .io_weight_win_33_ch2_33(conv_unit_1_io_weight_win_33_ch2_33),
    .io_weight_win_33_ch2_34(conv_unit_1_io_weight_win_33_ch2_34),
    .io_weight_win_33_ch2_35(conv_unit_1_io_weight_win_33_ch2_35),
    .io_weight_win_33_ch2_36(conv_unit_1_io_weight_win_33_ch2_36),
    .io_weight_win_33_ch2_37(conv_unit_1_io_weight_win_33_ch2_37),
    .io_weight_win_33_ch2_38(conv_unit_1_io_weight_win_33_ch2_38),
    .io_weight_win_33_ch2_39(conv_unit_1_io_weight_win_33_ch2_39),
    .io_weight_win_33_ch2_40(conv_unit_1_io_weight_win_33_ch2_40),
    .io_weight_win_33_ch2_41(conv_unit_1_io_weight_win_33_ch2_41),
    .io_weight_win_33_ch2_42(conv_unit_1_io_weight_win_33_ch2_42),
    .io_weight_win_33_ch2_43(conv_unit_1_io_weight_win_33_ch2_43),
    .io_weight_win_33_ch2_44(conv_unit_1_io_weight_win_33_ch2_44),
    .io_weight_win_33_ch2_45(conv_unit_1_io_weight_win_33_ch2_45),
    .io_weight_win_33_ch2_46(conv_unit_1_io_weight_win_33_ch2_46),
    .io_weight_win_33_ch2_47(conv_unit_1_io_weight_win_33_ch2_47),
    .io_weight_win_33_ch2_48(conv_unit_1_io_weight_win_33_ch2_48),
    .io_weight_win_33_ch2_49(conv_unit_1_io_weight_win_33_ch2_49),
    .io_weight_win_33_ch2_50(conv_unit_1_io_weight_win_33_ch2_50),
    .io_weight_win_33_ch2_51(conv_unit_1_io_weight_win_33_ch2_51),
    .io_weight_win_33_ch2_52(conv_unit_1_io_weight_win_33_ch2_52),
    .io_weight_win_33_ch2_53(conv_unit_1_io_weight_win_33_ch2_53),
    .io_weight_win_33_ch2_54(conv_unit_1_io_weight_win_33_ch2_54),
    .io_weight_win_33_ch2_55(conv_unit_1_io_weight_win_33_ch2_55),
    .io_weight_win_33_ch2_56(conv_unit_1_io_weight_win_33_ch2_56),
    .io_weight_win_33_ch2_57(conv_unit_1_io_weight_win_33_ch2_57),
    .io_weight_win_33_ch2_58(conv_unit_1_io_weight_win_33_ch2_58),
    .io_weight_win_33_ch2_59(conv_unit_1_io_weight_win_33_ch2_59),
    .io_weight_win_33_ch2_60(conv_unit_1_io_weight_win_33_ch2_60),
    .io_weight_win_33_ch2_61(conv_unit_1_io_weight_win_33_ch2_61),
    .io_weight_win_33_ch2_62(conv_unit_1_io_weight_win_33_ch2_62),
    .io_weight_win_33_ch2_63(conv_unit_1_io_weight_win_33_ch2_63),
    .io_weight_win_33_ch2_64(conv_unit_1_io_weight_win_33_ch2_64),
    .io_weight_win_33_ch2_65(conv_unit_1_io_weight_win_33_ch2_65),
    .io_weight_win_33_ch2_66(conv_unit_1_io_weight_win_33_ch2_66),
    .io_weight_win_33_ch2_67(conv_unit_1_io_weight_win_33_ch2_67),
    .io_weight_win_33_ch2_68(conv_unit_1_io_weight_win_33_ch2_68),
    .io_weight_win_33_ch2_69(conv_unit_1_io_weight_win_33_ch2_69),
    .io_weight_win_33_ch2_70(conv_unit_1_io_weight_win_33_ch2_70),
    .io_weight_win_33_ch2_71(conv_unit_1_io_weight_win_33_ch2_71),
    .io_bias1(conv_unit_1_io_bias1),
    .io_bias2(conv_unit_1_io_bias2),
    .io_bias_valid(conv_unit_1_io_bias_valid),
    .io_o_conv_ch1(conv_unit_1_io_o_conv_ch1),
    .io_o_conv_ch2(conv_unit_1_io_o_conv_ch2)
  );
  conv_unit conv_unit_2 ( // @[Conv.scala 18:47]
    .clock(conv_unit_2_clock),
    .io_ifm_win_33_0(conv_unit_2_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_unit_2_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_unit_2_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_unit_2_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_unit_2_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_unit_2_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_unit_2_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_unit_2_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_unit_2_io_ifm_win_33_8),
    .io_ifm_win_33_9(conv_unit_2_io_ifm_win_33_9),
    .io_ifm_win_33_10(conv_unit_2_io_ifm_win_33_10),
    .io_ifm_win_33_11(conv_unit_2_io_ifm_win_33_11),
    .io_ifm_win_33_12(conv_unit_2_io_ifm_win_33_12),
    .io_ifm_win_33_13(conv_unit_2_io_ifm_win_33_13),
    .io_ifm_win_33_14(conv_unit_2_io_ifm_win_33_14),
    .io_ifm_win_33_15(conv_unit_2_io_ifm_win_33_15),
    .io_ifm_win_33_16(conv_unit_2_io_ifm_win_33_16),
    .io_ifm_win_33_17(conv_unit_2_io_ifm_win_33_17),
    .io_ifm_win_33_18(conv_unit_2_io_ifm_win_33_18),
    .io_ifm_win_33_19(conv_unit_2_io_ifm_win_33_19),
    .io_ifm_win_33_20(conv_unit_2_io_ifm_win_33_20),
    .io_ifm_win_33_21(conv_unit_2_io_ifm_win_33_21),
    .io_ifm_win_33_22(conv_unit_2_io_ifm_win_33_22),
    .io_ifm_win_33_23(conv_unit_2_io_ifm_win_33_23),
    .io_ifm_win_33_24(conv_unit_2_io_ifm_win_33_24),
    .io_ifm_win_33_25(conv_unit_2_io_ifm_win_33_25),
    .io_ifm_win_33_26(conv_unit_2_io_ifm_win_33_26),
    .io_ifm_win_33_27(conv_unit_2_io_ifm_win_33_27),
    .io_ifm_win_33_28(conv_unit_2_io_ifm_win_33_28),
    .io_ifm_win_33_29(conv_unit_2_io_ifm_win_33_29),
    .io_ifm_win_33_30(conv_unit_2_io_ifm_win_33_30),
    .io_ifm_win_33_31(conv_unit_2_io_ifm_win_33_31),
    .io_ifm_win_33_32(conv_unit_2_io_ifm_win_33_32),
    .io_ifm_win_33_33(conv_unit_2_io_ifm_win_33_33),
    .io_ifm_win_33_34(conv_unit_2_io_ifm_win_33_34),
    .io_ifm_win_33_35(conv_unit_2_io_ifm_win_33_35),
    .io_ifm_win_33_36(conv_unit_2_io_ifm_win_33_36),
    .io_ifm_win_33_37(conv_unit_2_io_ifm_win_33_37),
    .io_ifm_win_33_38(conv_unit_2_io_ifm_win_33_38),
    .io_ifm_win_33_39(conv_unit_2_io_ifm_win_33_39),
    .io_ifm_win_33_40(conv_unit_2_io_ifm_win_33_40),
    .io_ifm_win_33_41(conv_unit_2_io_ifm_win_33_41),
    .io_ifm_win_33_42(conv_unit_2_io_ifm_win_33_42),
    .io_ifm_win_33_43(conv_unit_2_io_ifm_win_33_43),
    .io_ifm_win_33_44(conv_unit_2_io_ifm_win_33_44),
    .io_ifm_win_33_45(conv_unit_2_io_ifm_win_33_45),
    .io_ifm_win_33_46(conv_unit_2_io_ifm_win_33_46),
    .io_ifm_win_33_47(conv_unit_2_io_ifm_win_33_47),
    .io_ifm_win_33_48(conv_unit_2_io_ifm_win_33_48),
    .io_ifm_win_33_49(conv_unit_2_io_ifm_win_33_49),
    .io_ifm_win_33_50(conv_unit_2_io_ifm_win_33_50),
    .io_ifm_win_33_51(conv_unit_2_io_ifm_win_33_51),
    .io_ifm_win_33_52(conv_unit_2_io_ifm_win_33_52),
    .io_ifm_win_33_53(conv_unit_2_io_ifm_win_33_53),
    .io_ifm_win_33_54(conv_unit_2_io_ifm_win_33_54),
    .io_ifm_win_33_55(conv_unit_2_io_ifm_win_33_55),
    .io_ifm_win_33_56(conv_unit_2_io_ifm_win_33_56),
    .io_ifm_win_33_57(conv_unit_2_io_ifm_win_33_57),
    .io_ifm_win_33_58(conv_unit_2_io_ifm_win_33_58),
    .io_ifm_win_33_59(conv_unit_2_io_ifm_win_33_59),
    .io_ifm_win_33_60(conv_unit_2_io_ifm_win_33_60),
    .io_ifm_win_33_61(conv_unit_2_io_ifm_win_33_61),
    .io_ifm_win_33_62(conv_unit_2_io_ifm_win_33_62),
    .io_ifm_win_33_63(conv_unit_2_io_ifm_win_33_63),
    .io_ifm_win_33_64(conv_unit_2_io_ifm_win_33_64),
    .io_ifm_win_33_65(conv_unit_2_io_ifm_win_33_65),
    .io_ifm_win_33_66(conv_unit_2_io_ifm_win_33_66),
    .io_ifm_win_33_67(conv_unit_2_io_ifm_win_33_67),
    .io_ifm_win_33_68(conv_unit_2_io_ifm_win_33_68),
    .io_ifm_win_33_69(conv_unit_2_io_ifm_win_33_69),
    .io_ifm_win_33_70(conv_unit_2_io_ifm_win_33_70),
    .io_ifm_win_33_71(conv_unit_2_io_ifm_win_33_71),
    .io_weight_win_33_ch1_0(conv_unit_2_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_unit_2_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_unit_2_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_unit_2_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_unit_2_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_unit_2_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_unit_2_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_unit_2_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_unit_2_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch1_9(conv_unit_2_io_weight_win_33_ch1_9),
    .io_weight_win_33_ch1_10(conv_unit_2_io_weight_win_33_ch1_10),
    .io_weight_win_33_ch1_11(conv_unit_2_io_weight_win_33_ch1_11),
    .io_weight_win_33_ch1_12(conv_unit_2_io_weight_win_33_ch1_12),
    .io_weight_win_33_ch1_13(conv_unit_2_io_weight_win_33_ch1_13),
    .io_weight_win_33_ch1_14(conv_unit_2_io_weight_win_33_ch1_14),
    .io_weight_win_33_ch1_15(conv_unit_2_io_weight_win_33_ch1_15),
    .io_weight_win_33_ch1_16(conv_unit_2_io_weight_win_33_ch1_16),
    .io_weight_win_33_ch1_17(conv_unit_2_io_weight_win_33_ch1_17),
    .io_weight_win_33_ch1_18(conv_unit_2_io_weight_win_33_ch1_18),
    .io_weight_win_33_ch1_19(conv_unit_2_io_weight_win_33_ch1_19),
    .io_weight_win_33_ch1_20(conv_unit_2_io_weight_win_33_ch1_20),
    .io_weight_win_33_ch1_21(conv_unit_2_io_weight_win_33_ch1_21),
    .io_weight_win_33_ch1_22(conv_unit_2_io_weight_win_33_ch1_22),
    .io_weight_win_33_ch1_23(conv_unit_2_io_weight_win_33_ch1_23),
    .io_weight_win_33_ch1_24(conv_unit_2_io_weight_win_33_ch1_24),
    .io_weight_win_33_ch1_25(conv_unit_2_io_weight_win_33_ch1_25),
    .io_weight_win_33_ch1_26(conv_unit_2_io_weight_win_33_ch1_26),
    .io_weight_win_33_ch1_27(conv_unit_2_io_weight_win_33_ch1_27),
    .io_weight_win_33_ch1_28(conv_unit_2_io_weight_win_33_ch1_28),
    .io_weight_win_33_ch1_29(conv_unit_2_io_weight_win_33_ch1_29),
    .io_weight_win_33_ch1_30(conv_unit_2_io_weight_win_33_ch1_30),
    .io_weight_win_33_ch1_31(conv_unit_2_io_weight_win_33_ch1_31),
    .io_weight_win_33_ch1_32(conv_unit_2_io_weight_win_33_ch1_32),
    .io_weight_win_33_ch1_33(conv_unit_2_io_weight_win_33_ch1_33),
    .io_weight_win_33_ch1_34(conv_unit_2_io_weight_win_33_ch1_34),
    .io_weight_win_33_ch1_35(conv_unit_2_io_weight_win_33_ch1_35),
    .io_weight_win_33_ch1_36(conv_unit_2_io_weight_win_33_ch1_36),
    .io_weight_win_33_ch1_37(conv_unit_2_io_weight_win_33_ch1_37),
    .io_weight_win_33_ch1_38(conv_unit_2_io_weight_win_33_ch1_38),
    .io_weight_win_33_ch1_39(conv_unit_2_io_weight_win_33_ch1_39),
    .io_weight_win_33_ch1_40(conv_unit_2_io_weight_win_33_ch1_40),
    .io_weight_win_33_ch1_41(conv_unit_2_io_weight_win_33_ch1_41),
    .io_weight_win_33_ch1_42(conv_unit_2_io_weight_win_33_ch1_42),
    .io_weight_win_33_ch1_43(conv_unit_2_io_weight_win_33_ch1_43),
    .io_weight_win_33_ch1_44(conv_unit_2_io_weight_win_33_ch1_44),
    .io_weight_win_33_ch1_45(conv_unit_2_io_weight_win_33_ch1_45),
    .io_weight_win_33_ch1_46(conv_unit_2_io_weight_win_33_ch1_46),
    .io_weight_win_33_ch1_47(conv_unit_2_io_weight_win_33_ch1_47),
    .io_weight_win_33_ch1_48(conv_unit_2_io_weight_win_33_ch1_48),
    .io_weight_win_33_ch1_49(conv_unit_2_io_weight_win_33_ch1_49),
    .io_weight_win_33_ch1_50(conv_unit_2_io_weight_win_33_ch1_50),
    .io_weight_win_33_ch1_51(conv_unit_2_io_weight_win_33_ch1_51),
    .io_weight_win_33_ch1_52(conv_unit_2_io_weight_win_33_ch1_52),
    .io_weight_win_33_ch1_53(conv_unit_2_io_weight_win_33_ch1_53),
    .io_weight_win_33_ch1_54(conv_unit_2_io_weight_win_33_ch1_54),
    .io_weight_win_33_ch1_55(conv_unit_2_io_weight_win_33_ch1_55),
    .io_weight_win_33_ch1_56(conv_unit_2_io_weight_win_33_ch1_56),
    .io_weight_win_33_ch1_57(conv_unit_2_io_weight_win_33_ch1_57),
    .io_weight_win_33_ch1_58(conv_unit_2_io_weight_win_33_ch1_58),
    .io_weight_win_33_ch1_59(conv_unit_2_io_weight_win_33_ch1_59),
    .io_weight_win_33_ch1_60(conv_unit_2_io_weight_win_33_ch1_60),
    .io_weight_win_33_ch1_61(conv_unit_2_io_weight_win_33_ch1_61),
    .io_weight_win_33_ch1_62(conv_unit_2_io_weight_win_33_ch1_62),
    .io_weight_win_33_ch1_63(conv_unit_2_io_weight_win_33_ch1_63),
    .io_weight_win_33_ch1_64(conv_unit_2_io_weight_win_33_ch1_64),
    .io_weight_win_33_ch1_65(conv_unit_2_io_weight_win_33_ch1_65),
    .io_weight_win_33_ch1_66(conv_unit_2_io_weight_win_33_ch1_66),
    .io_weight_win_33_ch1_67(conv_unit_2_io_weight_win_33_ch1_67),
    .io_weight_win_33_ch1_68(conv_unit_2_io_weight_win_33_ch1_68),
    .io_weight_win_33_ch1_69(conv_unit_2_io_weight_win_33_ch1_69),
    .io_weight_win_33_ch1_70(conv_unit_2_io_weight_win_33_ch1_70),
    .io_weight_win_33_ch1_71(conv_unit_2_io_weight_win_33_ch1_71),
    .io_weight_win_33_ch2_0(conv_unit_2_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_unit_2_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_unit_2_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_unit_2_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_unit_2_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_unit_2_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_unit_2_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_unit_2_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_unit_2_io_weight_win_33_ch2_8),
    .io_weight_win_33_ch2_9(conv_unit_2_io_weight_win_33_ch2_9),
    .io_weight_win_33_ch2_10(conv_unit_2_io_weight_win_33_ch2_10),
    .io_weight_win_33_ch2_11(conv_unit_2_io_weight_win_33_ch2_11),
    .io_weight_win_33_ch2_12(conv_unit_2_io_weight_win_33_ch2_12),
    .io_weight_win_33_ch2_13(conv_unit_2_io_weight_win_33_ch2_13),
    .io_weight_win_33_ch2_14(conv_unit_2_io_weight_win_33_ch2_14),
    .io_weight_win_33_ch2_15(conv_unit_2_io_weight_win_33_ch2_15),
    .io_weight_win_33_ch2_16(conv_unit_2_io_weight_win_33_ch2_16),
    .io_weight_win_33_ch2_17(conv_unit_2_io_weight_win_33_ch2_17),
    .io_weight_win_33_ch2_18(conv_unit_2_io_weight_win_33_ch2_18),
    .io_weight_win_33_ch2_19(conv_unit_2_io_weight_win_33_ch2_19),
    .io_weight_win_33_ch2_20(conv_unit_2_io_weight_win_33_ch2_20),
    .io_weight_win_33_ch2_21(conv_unit_2_io_weight_win_33_ch2_21),
    .io_weight_win_33_ch2_22(conv_unit_2_io_weight_win_33_ch2_22),
    .io_weight_win_33_ch2_23(conv_unit_2_io_weight_win_33_ch2_23),
    .io_weight_win_33_ch2_24(conv_unit_2_io_weight_win_33_ch2_24),
    .io_weight_win_33_ch2_25(conv_unit_2_io_weight_win_33_ch2_25),
    .io_weight_win_33_ch2_26(conv_unit_2_io_weight_win_33_ch2_26),
    .io_weight_win_33_ch2_27(conv_unit_2_io_weight_win_33_ch2_27),
    .io_weight_win_33_ch2_28(conv_unit_2_io_weight_win_33_ch2_28),
    .io_weight_win_33_ch2_29(conv_unit_2_io_weight_win_33_ch2_29),
    .io_weight_win_33_ch2_30(conv_unit_2_io_weight_win_33_ch2_30),
    .io_weight_win_33_ch2_31(conv_unit_2_io_weight_win_33_ch2_31),
    .io_weight_win_33_ch2_32(conv_unit_2_io_weight_win_33_ch2_32),
    .io_weight_win_33_ch2_33(conv_unit_2_io_weight_win_33_ch2_33),
    .io_weight_win_33_ch2_34(conv_unit_2_io_weight_win_33_ch2_34),
    .io_weight_win_33_ch2_35(conv_unit_2_io_weight_win_33_ch2_35),
    .io_weight_win_33_ch2_36(conv_unit_2_io_weight_win_33_ch2_36),
    .io_weight_win_33_ch2_37(conv_unit_2_io_weight_win_33_ch2_37),
    .io_weight_win_33_ch2_38(conv_unit_2_io_weight_win_33_ch2_38),
    .io_weight_win_33_ch2_39(conv_unit_2_io_weight_win_33_ch2_39),
    .io_weight_win_33_ch2_40(conv_unit_2_io_weight_win_33_ch2_40),
    .io_weight_win_33_ch2_41(conv_unit_2_io_weight_win_33_ch2_41),
    .io_weight_win_33_ch2_42(conv_unit_2_io_weight_win_33_ch2_42),
    .io_weight_win_33_ch2_43(conv_unit_2_io_weight_win_33_ch2_43),
    .io_weight_win_33_ch2_44(conv_unit_2_io_weight_win_33_ch2_44),
    .io_weight_win_33_ch2_45(conv_unit_2_io_weight_win_33_ch2_45),
    .io_weight_win_33_ch2_46(conv_unit_2_io_weight_win_33_ch2_46),
    .io_weight_win_33_ch2_47(conv_unit_2_io_weight_win_33_ch2_47),
    .io_weight_win_33_ch2_48(conv_unit_2_io_weight_win_33_ch2_48),
    .io_weight_win_33_ch2_49(conv_unit_2_io_weight_win_33_ch2_49),
    .io_weight_win_33_ch2_50(conv_unit_2_io_weight_win_33_ch2_50),
    .io_weight_win_33_ch2_51(conv_unit_2_io_weight_win_33_ch2_51),
    .io_weight_win_33_ch2_52(conv_unit_2_io_weight_win_33_ch2_52),
    .io_weight_win_33_ch2_53(conv_unit_2_io_weight_win_33_ch2_53),
    .io_weight_win_33_ch2_54(conv_unit_2_io_weight_win_33_ch2_54),
    .io_weight_win_33_ch2_55(conv_unit_2_io_weight_win_33_ch2_55),
    .io_weight_win_33_ch2_56(conv_unit_2_io_weight_win_33_ch2_56),
    .io_weight_win_33_ch2_57(conv_unit_2_io_weight_win_33_ch2_57),
    .io_weight_win_33_ch2_58(conv_unit_2_io_weight_win_33_ch2_58),
    .io_weight_win_33_ch2_59(conv_unit_2_io_weight_win_33_ch2_59),
    .io_weight_win_33_ch2_60(conv_unit_2_io_weight_win_33_ch2_60),
    .io_weight_win_33_ch2_61(conv_unit_2_io_weight_win_33_ch2_61),
    .io_weight_win_33_ch2_62(conv_unit_2_io_weight_win_33_ch2_62),
    .io_weight_win_33_ch2_63(conv_unit_2_io_weight_win_33_ch2_63),
    .io_weight_win_33_ch2_64(conv_unit_2_io_weight_win_33_ch2_64),
    .io_weight_win_33_ch2_65(conv_unit_2_io_weight_win_33_ch2_65),
    .io_weight_win_33_ch2_66(conv_unit_2_io_weight_win_33_ch2_66),
    .io_weight_win_33_ch2_67(conv_unit_2_io_weight_win_33_ch2_67),
    .io_weight_win_33_ch2_68(conv_unit_2_io_weight_win_33_ch2_68),
    .io_weight_win_33_ch2_69(conv_unit_2_io_weight_win_33_ch2_69),
    .io_weight_win_33_ch2_70(conv_unit_2_io_weight_win_33_ch2_70),
    .io_weight_win_33_ch2_71(conv_unit_2_io_weight_win_33_ch2_71),
    .io_bias1(conv_unit_2_io_bias1),
    .io_bias2(conv_unit_2_io_bias2),
    .io_bias_valid(conv_unit_2_io_bias_valid),
    .io_o_conv_ch1(conv_unit_2_io_o_conv_ch1),
    .io_o_conv_ch2(conv_unit_2_io_o_conv_ch2)
  );
  conv_unit conv_unit_3 ( // @[Conv.scala 18:47]
    .clock(conv_unit_3_clock),
    .io_ifm_win_33_0(conv_unit_3_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_unit_3_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_unit_3_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_unit_3_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_unit_3_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_unit_3_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_unit_3_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_unit_3_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_unit_3_io_ifm_win_33_8),
    .io_ifm_win_33_9(conv_unit_3_io_ifm_win_33_9),
    .io_ifm_win_33_10(conv_unit_3_io_ifm_win_33_10),
    .io_ifm_win_33_11(conv_unit_3_io_ifm_win_33_11),
    .io_ifm_win_33_12(conv_unit_3_io_ifm_win_33_12),
    .io_ifm_win_33_13(conv_unit_3_io_ifm_win_33_13),
    .io_ifm_win_33_14(conv_unit_3_io_ifm_win_33_14),
    .io_ifm_win_33_15(conv_unit_3_io_ifm_win_33_15),
    .io_ifm_win_33_16(conv_unit_3_io_ifm_win_33_16),
    .io_ifm_win_33_17(conv_unit_3_io_ifm_win_33_17),
    .io_ifm_win_33_18(conv_unit_3_io_ifm_win_33_18),
    .io_ifm_win_33_19(conv_unit_3_io_ifm_win_33_19),
    .io_ifm_win_33_20(conv_unit_3_io_ifm_win_33_20),
    .io_ifm_win_33_21(conv_unit_3_io_ifm_win_33_21),
    .io_ifm_win_33_22(conv_unit_3_io_ifm_win_33_22),
    .io_ifm_win_33_23(conv_unit_3_io_ifm_win_33_23),
    .io_ifm_win_33_24(conv_unit_3_io_ifm_win_33_24),
    .io_ifm_win_33_25(conv_unit_3_io_ifm_win_33_25),
    .io_ifm_win_33_26(conv_unit_3_io_ifm_win_33_26),
    .io_ifm_win_33_27(conv_unit_3_io_ifm_win_33_27),
    .io_ifm_win_33_28(conv_unit_3_io_ifm_win_33_28),
    .io_ifm_win_33_29(conv_unit_3_io_ifm_win_33_29),
    .io_ifm_win_33_30(conv_unit_3_io_ifm_win_33_30),
    .io_ifm_win_33_31(conv_unit_3_io_ifm_win_33_31),
    .io_ifm_win_33_32(conv_unit_3_io_ifm_win_33_32),
    .io_ifm_win_33_33(conv_unit_3_io_ifm_win_33_33),
    .io_ifm_win_33_34(conv_unit_3_io_ifm_win_33_34),
    .io_ifm_win_33_35(conv_unit_3_io_ifm_win_33_35),
    .io_ifm_win_33_36(conv_unit_3_io_ifm_win_33_36),
    .io_ifm_win_33_37(conv_unit_3_io_ifm_win_33_37),
    .io_ifm_win_33_38(conv_unit_3_io_ifm_win_33_38),
    .io_ifm_win_33_39(conv_unit_3_io_ifm_win_33_39),
    .io_ifm_win_33_40(conv_unit_3_io_ifm_win_33_40),
    .io_ifm_win_33_41(conv_unit_3_io_ifm_win_33_41),
    .io_ifm_win_33_42(conv_unit_3_io_ifm_win_33_42),
    .io_ifm_win_33_43(conv_unit_3_io_ifm_win_33_43),
    .io_ifm_win_33_44(conv_unit_3_io_ifm_win_33_44),
    .io_ifm_win_33_45(conv_unit_3_io_ifm_win_33_45),
    .io_ifm_win_33_46(conv_unit_3_io_ifm_win_33_46),
    .io_ifm_win_33_47(conv_unit_3_io_ifm_win_33_47),
    .io_ifm_win_33_48(conv_unit_3_io_ifm_win_33_48),
    .io_ifm_win_33_49(conv_unit_3_io_ifm_win_33_49),
    .io_ifm_win_33_50(conv_unit_3_io_ifm_win_33_50),
    .io_ifm_win_33_51(conv_unit_3_io_ifm_win_33_51),
    .io_ifm_win_33_52(conv_unit_3_io_ifm_win_33_52),
    .io_ifm_win_33_53(conv_unit_3_io_ifm_win_33_53),
    .io_ifm_win_33_54(conv_unit_3_io_ifm_win_33_54),
    .io_ifm_win_33_55(conv_unit_3_io_ifm_win_33_55),
    .io_ifm_win_33_56(conv_unit_3_io_ifm_win_33_56),
    .io_ifm_win_33_57(conv_unit_3_io_ifm_win_33_57),
    .io_ifm_win_33_58(conv_unit_3_io_ifm_win_33_58),
    .io_ifm_win_33_59(conv_unit_3_io_ifm_win_33_59),
    .io_ifm_win_33_60(conv_unit_3_io_ifm_win_33_60),
    .io_ifm_win_33_61(conv_unit_3_io_ifm_win_33_61),
    .io_ifm_win_33_62(conv_unit_3_io_ifm_win_33_62),
    .io_ifm_win_33_63(conv_unit_3_io_ifm_win_33_63),
    .io_ifm_win_33_64(conv_unit_3_io_ifm_win_33_64),
    .io_ifm_win_33_65(conv_unit_3_io_ifm_win_33_65),
    .io_ifm_win_33_66(conv_unit_3_io_ifm_win_33_66),
    .io_ifm_win_33_67(conv_unit_3_io_ifm_win_33_67),
    .io_ifm_win_33_68(conv_unit_3_io_ifm_win_33_68),
    .io_ifm_win_33_69(conv_unit_3_io_ifm_win_33_69),
    .io_ifm_win_33_70(conv_unit_3_io_ifm_win_33_70),
    .io_ifm_win_33_71(conv_unit_3_io_ifm_win_33_71),
    .io_weight_win_33_ch1_0(conv_unit_3_io_weight_win_33_ch1_0),
    .io_weight_win_33_ch1_1(conv_unit_3_io_weight_win_33_ch1_1),
    .io_weight_win_33_ch1_2(conv_unit_3_io_weight_win_33_ch1_2),
    .io_weight_win_33_ch1_3(conv_unit_3_io_weight_win_33_ch1_3),
    .io_weight_win_33_ch1_4(conv_unit_3_io_weight_win_33_ch1_4),
    .io_weight_win_33_ch1_5(conv_unit_3_io_weight_win_33_ch1_5),
    .io_weight_win_33_ch1_6(conv_unit_3_io_weight_win_33_ch1_6),
    .io_weight_win_33_ch1_7(conv_unit_3_io_weight_win_33_ch1_7),
    .io_weight_win_33_ch1_8(conv_unit_3_io_weight_win_33_ch1_8),
    .io_weight_win_33_ch1_9(conv_unit_3_io_weight_win_33_ch1_9),
    .io_weight_win_33_ch1_10(conv_unit_3_io_weight_win_33_ch1_10),
    .io_weight_win_33_ch1_11(conv_unit_3_io_weight_win_33_ch1_11),
    .io_weight_win_33_ch1_12(conv_unit_3_io_weight_win_33_ch1_12),
    .io_weight_win_33_ch1_13(conv_unit_3_io_weight_win_33_ch1_13),
    .io_weight_win_33_ch1_14(conv_unit_3_io_weight_win_33_ch1_14),
    .io_weight_win_33_ch1_15(conv_unit_3_io_weight_win_33_ch1_15),
    .io_weight_win_33_ch1_16(conv_unit_3_io_weight_win_33_ch1_16),
    .io_weight_win_33_ch1_17(conv_unit_3_io_weight_win_33_ch1_17),
    .io_weight_win_33_ch1_18(conv_unit_3_io_weight_win_33_ch1_18),
    .io_weight_win_33_ch1_19(conv_unit_3_io_weight_win_33_ch1_19),
    .io_weight_win_33_ch1_20(conv_unit_3_io_weight_win_33_ch1_20),
    .io_weight_win_33_ch1_21(conv_unit_3_io_weight_win_33_ch1_21),
    .io_weight_win_33_ch1_22(conv_unit_3_io_weight_win_33_ch1_22),
    .io_weight_win_33_ch1_23(conv_unit_3_io_weight_win_33_ch1_23),
    .io_weight_win_33_ch1_24(conv_unit_3_io_weight_win_33_ch1_24),
    .io_weight_win_33_ch1_25(conv_unit_3_io_weight_win_33_ch1_25),
    .io_weight_win_33_ch1_26(conv_unit_3_io_weight_win_33_ch1_26),
    .io_weight_win_33_ch1_27(conv_unit_3_io_weight_win_33_ch1_27),
    .io_weight_win_33_ch1_28(conv_unit_3_io_weight_win_33_ch1_28),
    .io_weight_win_33_ch1_29(conv_unit_3_io_weight_win_33_ch1_29),
    .io_weight_win_33_ch1_30(conv_unit_3_io_weight_win_33_ch1_30),
    .io_weight_win_33_ch1_31(conv_unit_3_io_weight_win_33_ch1_31),
    .io_weight_win_33_ch1_32(conv_unit_3_io_weight_win_33_ch1_32),
    .io_weight_win_33_ch1_33(conv_unit_3_io_weight_win_33_ch1_33),
    .io_weight_win_33_ch1_34(conv_unit_3_io_weight_win_33_ch1_34),
    .io_weight_win_33_ch1_35(conv_unit_3_io_weight_win_33_ch1_35),
    .io_weight_win_33_ch1_36(conv_unit_3_io_weight_win_33_ch1_36),
    .io_weight_win_33_ch1_37(conv_unit_3_io_weight_win_33_ch1_37),
    .io_weight_win_33_ch1_38(conv_unit_3_io_weight_win_33_ch1_38),
    .io_weight_win_33_ch1_39(conv_unit_3_io_weight_win_33_ch1_39),
    .io_weight_win_33_ch1_40(conv_unit_3_io_weight_win_33_ch1_40),
    .io_weight_win_33_ch1_41(conv_unit_3_io_weight_win_33_ch1_41),
    .io_weight_win_33_ch1_42(conv_unit_3_io_weight_win_33_ch1_42),
    .io_weight_win_33_ch1_43(conv_unit_3_io_weight_win_33_ch1_43),
    .io_weight_win_33_ch1_44(conv_unit_3_io_weight_win_33_ch1_44),
    .io_weight_win_33_ch1_45(conv_unit_3_io_weight_win_33_ch1_45),
    .io_weight_win_33_ch1_46(conv_unit_3_io_weight_win_33_ch1_46),
    .io_weight_win_33_ch1_47(conv_unit_3_io_weight_win_33_ch1_47),
    .io_weight_win_33_ch1_48(conv_unit_3_io_weight_win_33_ch1_48),
    .io_weight_win_33_ch1_49(conv_unit_3_io_weight_win_33_ch1_49),
    .io_weight_win_33_ch1_50(conv_unit_3_io_weight_win_33_ch1_50),
    .io_weight_win_33_ch1_51(conv_unit_3_io_weight_win_33_ch1_51),
    .io_weight_win_33_ch1_52(conv_unit_3_io_weight_win_33_ch1_52),
    .io_weight_win_33_ch1_53(conv_unit_3_io_weight_win_33_ch1_53),
    .io_weight_win_33_ch1_54(conv_unit_3_io_weight_win_33_ch1_54),
    .io_weight_win_33_ch1_55(conv_unit_3_io_weight_win_33_ch1_55),
    .io_weight_win_33_ch1_56(conv_unit_3_io_weight_win_33_ch1_56),
    .io_weight_win_33_ch1_57(conv_unit_3_io_weight_win_33_ch1_57),
    .io_weight_win_33_ch1_58(conv_unit_3_io_weight_win_33_ch1_58),
    .io_weight_win_33_ch1_59(conv_unit_3_io_weight_win_33_ch1_59),
    .io_weight_win_33_ch1_60(conv_unit_3_io_weight_win_33_ch1_60),
    .io_weight_win_33_ch1_61(conv_unit_3_io_weight_win_33_ch1_61),
    .io_weight_win_33_ch1_62(conv_unit_3_io_weight_win_33_ch1_62),
    .io_weight_win_33_ch1_63(conv_unit_3_io_weight_win_33_ch1_63),
    .io_weight_win_33_ch1_64(conv_unit_3_io_weight_win_33_ch1_64),
    .io_weight_win_33_ch1_65(conv_unit_3_io_weight_win_33_ch1_65),
    .io_weight_win_33_ch1_66(conv_unit_3_io_weight_win_33_ch1_66),
    .io_weight_win_33_ch1_67(conv_unit_3_io_weight_win_33_ch1_67),
    .io_weight_win_33_ch1_68(conv_unit_3_io_weight_win_33_ch1_68),
    .io_weight_win_33_ch1_69(conv_unit_3_io_weight_win_33_ch1_69),
    .io_weight_win_33_ch1_70(conv_unit_3_io_weight_win_33_ch1_70),
    .io_weight_win_33_ch1_71(conv_unit_3_io_weight_win_33_ch1_71),
    .io_weight_win_33_ch2_0(conv_unit_3_io_weight_win_33_ch2_0),
    .io_weight_win_33_ch2_1(conv_unit_3_io_weight_win_33_ch2_1),
    .io_weight_win_33_ch2_2(conv_unit_3_io_weight_win_33_ch2_2),
    .io_weight_win_33_ch2_3(conv_unit_3_io_weight_win_33_ch2_3),
    .io_weight_win_33_ch2_4(conv_unit_3_io_weight_win_33_ch2_4),
    .io_weight_win_33_ch2_5(conv_unit_3_io_weight_win_33_ch2_5),
    .io_weight_win_33_ch2_6(conv_unit_3_io_weight_win_33_ch2_6),
    .io_weight_win_33_ch2_7(conv_unit_3_io_weight_win_33_ch2_7),
    .io_weight_win_33_ch2_8(conv_unit_3_io_weight_win_33_ch2_8),
    .io_weight_win_33_ch2_9(conv_unit_3_io_weight_win_33_ch2_9),
    .io_weight_win_33_ch2_10(conv_unit_3_io_weight_win_33_ch2_10),
    .io_weight_win_33_ch2_11(conv_unit_3_io_weight_win_33_ch2_11),
    .io_weight_win_33_ch2_12(conv_unit_3_io_weight_win_33_ch2_12),
    .io_weight_win_33_ch2_13(conv_unit_3_io_weight_win_33_ch2_13),
    .io_weight_win_33_ch2_14(conv_unit_3_io_weight_win_33_ch2_14),
    .io_weight_win_33_ch2_15(conv_unit_3_io_weight_win_33_ch2_15),
    .io_weight_win_33_ch2_16(conv_unit_3_io_weight_win_33_ch2_16),
    .io_weight_win_33_ch2_17(conv_unit_3_io_weight_win_33_ch2_17),
    .io_weight_win_33_ch2_18(conv_unit_3_io_weight_win_33_ch2_18),
    .io_weight_win_33_ch2_19(conv_unit_3_io_weight_win_33_ch2_19),
    .io_weight_win_33_ch2_20(conv_unit_3_io_weight_win_33_ch2_20),
    .io_weight_win_33_ch2_21(conv_unit_3_io_weight_win_33_ch2_21),
    .io_weight_win_33_ch2_22(conv_unit_3_io_weight_win_33_ch2_22),
    .io_weight_win_33_ch2_23(conv_unit_3_io_weight_win_33_ch2_23),
    .io_weight_win_33_ch2_24(conv_unit_3_io_weight_win_33_ch2_24),
    .io_weight_win_33_ch2_25(conv_unit_3_io_weight_win_33_ch2_25),
    .io_weight_win_33_ch2_26(conv_unit_3_io_weight_win_33_ch2_26),
    .io_weight_win_33_ch2_27(conv_unit_3_io_weight_win_33_ch2_27),
    .io_weight_win_33_ch2_28(conv_unit_3_io_weight_win_33_ch2_28),
    .io_weight_win_33_ch2_29(conv_unit_3_io_weight_win_33_ch2_29),
    .io_weight_win_33_ch2_30(conv_unit_3_io_weight_win_33_ch2_30),
    .io_weight_win_33_ch2_31(conv_unit_3_io_weight_win_33_ch2_31),
    .io_weight_win_33_ch2_32(conv_unit_3_io_weight_win_33_ch2_32),
    .io_weight_win_33_ch2_33(conv_unit_3_io_weight_win_33_ch2_33),
    .io_weight_win_33_ch2_34(conv_unit_3_io_weight_win_33_ch2_34),
    .io_weight_win_33_ch2_35(conv_unit_3_io_weight_win_33_ch2_35),
    .io_weight_win_33_ch2_36(conv_unit_3_io_weight_win_33_ch2_36),
    .io_weight_win_33_ch2_37(conv_unit_3_io_weight_win_33_ch2_37),
    .io_weight_win_33_ch2_38(conv_unit_3_io_weight_win_33_ch2_38),
    .io_weight_win_33_ch2_39(conv_unit_3_io_weight_win_33_ch2_39),
    .io_weight_win_33_ch2_40(conv_unit_3_io_weight_win_33_ch2_40),
    .io_weight_win_33_ch2_41(conv_unit_3_io_weight_win_33_ch2_41),
    .io_weight_win_33_ch2_42(conv_unit_3_io_weight_win_33_ch2_42),
    .io_weight_win_33_ch2_43(conv_unit_3_io_weight_win_33_ch2_43),
    .io_weight_win_33_ch2_44(conv_unit_3_io_weight_win_33_ch2_44),
    .io_weight_win_33_ch2_45(conv_unit_3_io_weight_win_33_ch2_45),
    .io_weight_win_33_ch2_46(conv_unit_3_io_weight_win_33_ch2_46),
    .io_weight_win_33_ch2_47(conv_unit_3_io_weight_win_33_ch2_47),
    .io_weight_win_33_ch2_48(conv_unit_3_io_weight_win_33_ch2_48),
    .io_weight_win_33_ch2_49(conv_unit_3_io_weight_win_33_ch2_49),
    .io_weight_win_33_ch2_50(conv_unit_3_io_weight_win_33_ch2_50),
    .io_weight_win_33_ch2_51(conv_unit_3_io_weight_win_33_ch2_51),
    .io_weight_win_33_ch2_52(conv_unit_3_io_weight_win_33_ch2_52),
    .io_weight_win_33_ch2_53(conv_unit_3_io_weight_win_33_ch2_53),
    .io_weight_win_33_ch2_54(conv_unit_3_io_weight_win_33_ch2_54),
    .io_weight_win_33_ch2_55(conv_unit_3_io_weight_win_33_ch2_55),
    .io_weight_win_33_ch2_56(conv_unit_3_io_weight_win_33_ch2_56),
    .io_weight_win_33_ch2_57(conv_unit_3_io_weight_win_33_ch2_57),
    .io_weight_win_33_ch2_58(conv_unit_3_io_weight_win_33_ch2_58),
    .io_weight_win_33_ch2_59(conv_unit_3_io_weight_win_33_ch2_59),
    .io_weight_win_33_ch2_60(conv_unit_3_io_weight_win_33_ch2_60),
    .io_weight_win_33_ch2_61(conv_unit_3_io_weight_win_33_ch2_61),
    .io_weight_win_33_ch2_62(conv_unit_3_io_weight_win_33_ch2_62),
    .io_weight_win_33_ch2_63(conv_unit_3_io_weight_win_33_ch2_63),
    .io_weight_win_33_ch2_64(conv_unit_3_io_weight_win_33_ch2_64),
    .io_weight_win_33_ch2_65(conv_unit_3_io_weight_win_33_ch2_65),
    .io_weight_win_33_ch2_66(conv_unit_3_io_weight_win_33_ch2_66),
    .io_weight_win_33_ch2_67(conv_unit_3_io_weight_win_33_ch2_67),
    .io_weight_win_33_ch2_68(conv_unit_3_io_weight_win_33_ch2_68),
    .io_weight_win_33_ch2_69(conv_unit_3_io_weight_win_33_ch2_69),
    .io_weight_win_33_ch2_70(conv_unit_3_io_weight_win_33_ch2_70),
    .io_weight_win_33_ch2_71(conv_unit_3_io_weight_win_33_ch2_71),
    .io_bias1(conv_unit_3_io_bias1),
    .io_bias2(conv_unit_3_io_bias2),
    .io_bias_valid(conv_unit_3_io_bias_valid),
    .io_o_conv_ch1(conv_unit_3_io_o_conv_ch1),
    .io_o_conv_ch2(conv_unit_3_io_o_conv_ch2)
  );
  assign io_conv_o_0 = conv_unit_0_io_o_conv_ch1; // @[Conv.scala 28:26]
  assign io_conv_o_1 = conv_unit_0_io_o_conv_ch2; // @[Conv.scala 29:30]
  assign io_conv_o_2 = conv_unit_1_io_o_conv_ch1; // @[Conv.scala 28:26]
  assign io_conv_o_3 = conv_unit_1_io_o_conv_ch2; // @[Conv.scala 29:30]
  assign io_conv_o_4 = conv_unit_2_io_o_conv_ch1; // @[Conv.scala 28:26]
  assign io_conv_o_5 = conv_unit_2_io_o_conv_ch2; // @[Conv.scala 29:30]
  assign io_conv_o_6 = conv_unit_3_io_o_conv_ch1; // @[Conv.scala 28:26]
  assign io_conv_o_7 = conv_unit_3_io_o_conv_ch2; // @[Conv.scala 29:30]
  assign conv_unit_0_clock = clock;
  assign conv_unit_0_io_ifm_win_33_0 = io_ifm_win_33_0; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_1 = io_ifm_win_33_1; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_2 = io_ifm_win_33_2; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_3 = io_ifm_win_33_3; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_4 = io_ifm_win_33_4; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_5 = io_ifm_win_33_5; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_6 = io_ifm_win_33_6; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_7 = io_ifm_win_33_7; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_8 = io_ifm_win_33_8; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_9 = io_ifm_win_33_9; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_10 = io_ifm_win_33_10; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_11 = io_ifm_win_33_11; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_12 = io_ifm_win_33_12; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_13 = io_ifm_win_33_13; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_14 = io_ifm_win_33_14; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_15 = io_ifm_win_33_15; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_16 = io_ifm_win_33_16; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_17 = io_ifm_win_33_17; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_18 = io_ifm_win_33_18; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_19 = io_ifm_win_33_19; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_20 = io_ifm_win_33_20; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_21 = io_ifm_win_33_21; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_22 = io_ifm_win_33_22; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_23 = io_ifm_win_33_23; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_24 = io_ifm_win_33_24; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_25 = io_ifm_win_33_25; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_26 = io_ifm_win_33_26; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_27 = io_ifm_win_33_27; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_28 = io_ifm_win_33_28; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_29 = io_ifm_win_33_29; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_30 = io_ifm_win_33_30; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_31 = io_ifm_win_33_31; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_32 = io_ifm_win_33_32; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_33 = io_ifm_win_33_33; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_34 = io_ifm_win_33_34; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_35 = io_ifm_win_33_35; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_36 = io_ifm_win_33_36; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_37 = io_ifm_win_33_37; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_38 = io_ifm_win_33_38; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_39 = io_ifm_win_33_39; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_40 = io_ifm_win_33_40; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_41 = io_ifm_win_33_41; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_42 = io_ifm_win_33_42; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_43 = io_ifm_win_33_43; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_44 = io_ifm_win_33_44; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_45 = io_ifm_win_33_45; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_46 = io_ifm_win_33_46; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_47 = io_ifm_win_33_47; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_48 = io_ifm_win_33_48; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_49 = io_ifm_win_33_49; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_50 = io_ifm_win_33_50; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_51 = io_ifm_win_33_51; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_52 = io_ifm_win_33_52; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_53 = io_ifm_win_33_53; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_54 = io_ifm_win_33_54; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_55 = io_ifm_win_33_55; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_56 = io_ifm_win_33_56; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_57 = io_ifm_win_33_57; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_58 = io_ifm_win_33_58; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_59 = io_ifm_win_33_59; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_60 = io_ifm_win_33_60; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_61 = io_ifm_win_33_61; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_62 = io_ifm_win_33_62; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_63 = io_ifm_win_33_63; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_64 = io_ifm_win_33_64; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_65 = io_ifm_win_33_65; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_66 = io_ifm_win_33_66; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_67 = io_ifm_win_33_67; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_68 = io_ifm_win_33_68; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_69 = io_ifm_win_33_69; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_70 = io_ifm_win_33_70; // @[Conv.scala 20:36]
  assign conv_unit_0_io_ifm_win_33_71 = io_ifm_win_33_71; // @[Conv.scala 20:36]
  assign conv_unit_0_io_weight_win_33_ch1_0 = io_weight_win_33_0; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_1 = io_weight_win_33_1; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_2 = io_weight_win_33_2; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_3 = io_weight_win_33_3; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_4 = io_weight_win_33_4; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_5 = io_weight_win_33_5; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_6 = io_weight_win_33_6; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_7 = io_weight_win_33_7; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_8 = io_weight_win_33_8; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_9 = io_weight_win_33_9; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_10 = io_weight_win_33_10; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_11 = io_weight_win_33_11; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_12 = io_weight_win_33_12; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_13 = io_weight_win_33_13; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_14 = io_weight_win_33_14; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_15 = io_weight_win_33_15; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_16 = io_weight_win_33_16; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_17 = io_weight_win_33_17; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_18 = io_weight_win_33_18; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_19 = io_weight_win_33_19; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_20 = io_weight_win_33_20; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_21 = io_weight_win_33_21; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_22 = io_weight_win_33_22; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_23 = io_weight_win_33_23; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_24 = io_weight_win_33_24; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_25 = io_weight_win_33_25; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_26 = io_weight_win_33_26; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_27 = io_weight_win_33_27; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_28 = io_weight_win_33_28; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_29 = io_weight_win_33_29; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_30 = io_weight_win_33_30; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_31 = io_weight_win_33_31; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_32 = io_weight_win_33_32; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_33 = io_weight_win_33_33; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_34 = io_weight_win_33_34; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_35 = io_weight_win_33_35; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_36 = io_weight_win_33_36; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_37 = io_weight_win_33_37; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_38 = io_weight_win_33_38; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_39 = io_weight_win_33_39; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_40 = io_weight_win_33_40; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_41 = io_weight_win_33_41; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_42 = io_weight_win_33_42; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_43 = io_weight_win_33_43; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_44 = io_weight_win_33_44; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_45 = io_weight_win_33_45; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_46 = io_weight_win_33_46; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_47 = io_weight_win_33_47; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_48 = io_weight_win_33_48; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_49 = io_weight_win_33_49; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_50 = io_weight_win_33_50; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_51 = io_weight_win_33_51; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_52 = io_weight_win_33_52; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_53 = io_weight_win_33_53; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_54 = io_weight_win_33_54; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_55 = io_weight_win_33_55; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_56 = io_weight_win_33_56; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_57 = io_weight_win_33_57; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_58 = io_weight_win_33_58; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_59 = io_weight_win_33_59; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_60 = io_weight_win_33_60; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_61 = io_weight_win_33_61; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_62 = io_weight_win_33_62; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_63 = io_weight_win_33_63; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_64 = io_weight_win_33_64; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_65 = io_weight_win_33_65; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_66 = io_weight_win_33_66; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_67 = io_weight_win_33_67; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_68 = io_weight_win_33_68; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_69 = io_weight_win_33_69; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_70 = io_weight_win_33_70; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch1_71 = io_weight_win_33_71; // @[Conv.scala 22:50]
  assign conv_unit_0_io_weight_win_33_ch2_0 = io_weight_win_33_72; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_1 = io_weight_win_33_73; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_2 = io_weight_win_33_74; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_3 = io_weight_win_33_75; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_4 = io_weight_win_33_76; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_5 = io_weight_win_33_77; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_6 = io_weight_win_33_78; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_7 = io_weight_win_33_79; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_8 = io_weight_win_33_80; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_9 = io_weight_win_33_81; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_10 = io_weight_win_33_82; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_11 = io_weight_win_33_83; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_12 = io_weight_win_33_84; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_13 = io_weight_win_33_85; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_14 = io_weight_win_33_86; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_15 = io_weight_win_33_87; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_16 = io_weight_win_33_88; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_17 = io_weight_win_33_89; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_18 = io_weight_win_33_90; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_19 = io_weight_win_33_91; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_20 = io_weight_win_33_92; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_21 = io_weight_win_33_93; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_22 = io_weight_win_33_94; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_23 = io_weight_win_33_95; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_24 = io_weight_win_33_96; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_25 = io_weight_win_33_97; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_26 = io_weight_win_33_98; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_27 = io_weight_win_33_99; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_28 = io_weight_win_33_100; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_29 = io_weight_win_33_101; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_30 = io_weight_win_33_102; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_31 = io_weight_win_33_103; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_32 = io_weight_win_33_104; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_33 = io_weight_win_33_105; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_34 = io_weight_win_33_106; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_35 = io_weight_win_33_107; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_36 = io_weight_win_33_108; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_37 = io_weight_win_33_109; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_38 = io_weight_win_33_110; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_39 = io_weight_win_33_111; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_40 = io_weight_win_33_112; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_41 = io_weight_win_33_113; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_42 = io_weight_win_33_114; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_43 = io_weight_win_33_115; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_44 = io_weight_win_33_116; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_45 = io_weight_win_33_117; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_46 = io_weight_win_33_118; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_47 = io_weight_win_33_119; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_48 = io_weight_win_33_120; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_49 = io_weight_win_33_121; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_50 = io_weight_win_33_122; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_51 = io_weight_win_33_123; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_52 = io_weight_win_33_124; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_53 = io_weight_win_33_125; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_54 = io_weight_win_33_126; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_55 = io_weight_win_33_127; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_56 = io_weight_win_33_128; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_57 = io_weight_win_33_129; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_58 = io_weight_win_33_130; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_59 = io_weight_win_33_131; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_60 = io_weight_win_33_132; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_61 = io_weight_win_33_133; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_62 = io_weight_win_33_134; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_63 = io_weight_win_33_135; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_64 = io_weight_win_33_136; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_65 = io_weight_win_33_137; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_66 = io_weight_win_33_138; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_67 = io_weight_win_33_139; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_68 = io_weight_win_33_140; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_69 = io_weight_win_33_141; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_70 = io_weight_win_33_142; // @[Conv.scala 23:50]
  assign conv_unit_0_io_weight_win_33_ch2_71 = io_weight_win_33_143; // @[Conv.scala 23:50]
  assign conv_unit_0_io_bias1 = io_bias_data_0; // @[Conv.scala 25:31]
  assign conv_unit_0_io_bias2 = io_bias_data_1; // @[Conv.scala 26:31]
  assign conv_unit_0_io_bias_valid = io_bias_valid; // @[Conv.scala 27:36]
  assign conv_unit_1_clock = clock;
  assign conv_unit_1_io_ifm_win_33_0 = io_ifm_win_33_0; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_1 = io_ifm_win_33_1; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_2 = io_ifm_win_33_2; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_3 = io_ifm_win_33_3; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_4 = io_ifm_win_33_4; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_5 = io_ifm_win_33_5; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_6 = io_ifm_win_33_6; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_7 = io_ifm_win_33_7; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_8 = io_ifm_win_33_8; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_9 = io_ifm_win_33_9; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_10 = io_ifm_win_33_10; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_11 = io_ifm_win_33_11; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_12 = io_ifm_win_33_12; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_13 = io_ifm_win_33_13; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_14 = io_ifm_win_33_14; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_15 = io_ifm_win_33_15; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_16 = io_ifm_win_33_16; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_17 = io_ifm_win_33_17; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_18 = io_ifm_win_33_18; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_19 = io_ifm_win_33_19; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_20 = io_ifm_win_33_20; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_21 = io_ifm_win_33_21; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_22 = io_ifm_win_33_22; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_23 = io_ifm_win_33_23; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_24 = io_ifm_win_33_24; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_25 = io_ifm_win_33_25; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_26 = io_ifm_win_33_26; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_27 = io_ifm_win_33_27; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_28 = io_ifm_win_33_28; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_29 = io_ifm_win_33_29; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_30 = io_ifm_win_33_30; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_31 = io_ifm_win_33_31; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_32 = io_ifm_win_33_32; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_33 = io_ifm_win_33_33; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_34 = io_ifm_win_33_34; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_35 = io_ifm_win_33_35; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_36 = io_ifm_win_33_36; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_37 = io_ifm_win_33_37; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_38 = io_ifm_win_33_38; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_39 = io_ifm_win_33_39; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_40 = io_ifm_win_33_40; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_41 = io_ifm_win_33_41; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_42 = io_ifm_win_33_42; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_43 = io_ifm_win_33_43; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_44 = io_ifm_win_33_44; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_45 = io_ifm_win_33_45; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_46 = io_ifm_win_33_46; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_47 = io_ifm_win_33_47; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_48 = io_ifm_win_33_48; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_49 = io_ifm_win_33_49; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_50 = io_ifm_win_33_50; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_51 = io_ifm_win_33_51; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_52 = io_ifm_win_33_52; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_53 = io_ifm_win_33_53; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_54 = io_ifm_win_33_54; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_55 = io_ifm_win_33_55; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_56 = io_ifm_win_33_56; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_57 = io_ifm_win_33_57; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_58 = io_ifm_win_33_58; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_59 = io_ifm_win_33_59; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_60 = io_ifm_win_33_60; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_61 = io_ifm_win_33_61; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_62 = io_ifm_win_33_62; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_63 = io_ifm_win_33_63; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_64 = io_ifm_win_33_64; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_65 = io_ifm_win_33_65; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_66 = io_ifm_win_33_66; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_67 = io_ifm_win_33_67; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_68 = io_ifm_win_33_68; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_69 = io_ifm_win_33_69; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_70 = io_ifm_win_33_70; // @[Conv.scala 20:36]
  assign conv_unit_1_io_ifm_win_33_71 = io_ifm_win_33_71; // @[Conv.scala 20:36]
  assign conv_unit_1_io_weight_win_33_ch1_0 = io_weight_win_33_144; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_1 = io_weight_win_33_145; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_2 = io_weight_win_33_146; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_3 = io_weight_win_33_147; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_4 = io_weight_win_33_148; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_5 = io_weight_win_33_149; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_6 = io_weight_win_33_150; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_7 = io_weight_win_33_151; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_8 = io_weight_win_33_152; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_9 = io_weight_win_33_153; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_10 = io_weight_win_33_154; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_11 = io_weight_win_33_155; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_12 = io_weight_win_33_156; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_13 = io_weight_win_33_157; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_14 = io_weight_win_33_158; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_15 = io_weight_win_33_159; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_16 = io_weight_win_33_160; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_17 = io_weight_win_33_161; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_18 = io_weight_win_33_162; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_19 = io_weight_win_33_163; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_20 = io_weight_win_33_164; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_21 = io_weight_win_33_165; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_22 = io_weight_win_33_166; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_23 = io_weight_win_33_167; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_24 = io_weight_win_33_168; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_25 = io_weight_win_33_169; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_26 = io_weight_win_33_170; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_27 = io_weight_win_33_171; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_28 = io_weight_win_33_172; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_29 = io_weight_win_33_173; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_30 = io_weight_win_33_174; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_31 = io_weight_win_33_175; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_32 = io_weight_win_33_176; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_33 = io_weight_win_33_177; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_34 = io_weight_win_33_178; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_35 = io_weight_win_33_179; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_36 = io_weight_win_33_180; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_37 = io_weight_win_33_181; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_38 = io_weight_win_33_182; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_39 = io_weight_win_33_183; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_40 = io_weight_win_33_184; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_41 = io_weight_win_33_185; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_42 = io_weight_win_33_186; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_43 = io_weight_win_33_187; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_44 = io_weight_win_33_188; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_45 = io_weight_win_33_189; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_46 = io_weight_win_33_190; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_47 = io_weight_win_33_191; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_48 = io_weight_win_33_192; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_49 = io_weight_win_33_193; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_50 = io_weight_win_33_194; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_51 = io_weight_win_33_195; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_52 = io_weight_win_33_196; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_53 = io_weight_win_33_197; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_54 = io_weight_win_33_198; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_55 = io_weight_win_33_199; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_56 = io_weight_win_33_200; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_57 = io_weight_win_33_201; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_58 = io_weight_win_33_202; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_59 = io_weight_win_33_203; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_60 = io_weight_win_33_204; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_61 = io_weight_win_33_205; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_62 = io_weight_win_33_206; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_63 = io_weight_win_33_207; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_64 = io_weight_win_33_208; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_65 = io_weight_win_33_209; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_66 = io_weight_win_33_210; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_67 = io_weight_win_33_211; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_68 = io_weight_win_33_212; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_69 = io_weight_win_33_213; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_70 = io_weight_win_33_214; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch1_71 = io_weight_win_33_215; // @[Conv.scala 22:50]
  assign conv_unit_1_io_weight_win_33_ch2_0 = io_weight_win_33_216; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_1 = io_weight_win_33_217; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_2 = io_weight_win_33_218; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_3 = io_weight_win_33_219; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_4 = io_weight_win_33_220; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_5 = io_weight_win_33_221; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_6 = io_weight_win_33_222; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_7 = io_weight_win_33_223; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_8 = io_weight_win_33_224; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_9 = io_weight_win_33_225; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_10 = io_weight_win_33_226; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_11 = io_weight_win_33_227; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_12 = io_weight_win_33_228; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_13 = io_weight_win_33_229; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_14 = io_weight_win_33_230; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_15 = io_weight_win_33_231; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_16 = io_weight_win_33_232; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_17 = io_weight_win_33_233; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_18 = io_weight_win_33_234; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_19 = io_weight_win_33_235; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_20 = io_weight_win_33_236; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_21 = io_weight_win_33_237; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_22 = io_weight_win_33_238; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_23 = io_weight_win_33_239; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_24 = io_weight_win_33_240; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_25 = io_weight_win_33_241; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_26 = io_weight_win_33_242; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_27 = io_weight_win_33_243; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_28 = io_weight_win_33_244; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_29 = io_weight_win_33_245; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_30 = io_weight_win_33_246; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_31 = io_weight_win_33_247; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_32 = io_weight_win_33_248; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_33 = io_weight_win_33_249; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_34 = io_weight_win_33_250; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_35 = io_weight_win_33_251; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_36 = io_weight_win_33_252; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_37 = io_weight_win_33_253; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_38 = io_weight_win_33_254; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_39 = io_weight_win_33_255; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_40 = io_weight_win_33_256; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_41 = io_weight_win_33_257; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_42 = io_weight_win_33_258; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_43 = io_weight_win_33_259; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_44 = io_weight_win_33_260; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_45 = io_weight_win_33_261; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_46 = io_weight_win_33_262; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_47 = io_weight_win_33_263; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_48 = io_weight_win_33_264; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_49 = io_weight_win_33_265; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_50 = io_weight_win_33_266; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_51 = io_weight_win_33_267; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_52 = io_weight_win_33_268; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_53 = io_weight_win_33_269; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_54 = io_weight_win_33_270; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_55 = io_weight_win_33_271; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_56 = io_weight_win_33_272; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_57 = io_weight_win_33_273; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_58 = io_weight_win_33_274; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_59 = io_weight_win_33_275; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_60 = io_weight_win_33_276; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_61 = io_weight_win_33_277; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_62 = io_weight_win_33_278; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_63 = io_weight_win_33_279; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_64 = io_weight_win_33_280; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_65 = io_weight_win_33_281; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_66 = io_weight_win_33_282; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_67 = io_weight_win_33_283; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_68 = io_weight_win_33_284; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_69 = io_weight_win_33_285; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_70 = io_weight_win_33_286; // @[Conv.scala 23:50]
  assign conv_unit_1_io_weight_win_33_ch2_71 = io_weight_win_33_287; // @[Conv.scala 23:50]
  assign conv_unit_1_io_bias1 = io_bias_data_2; // @[Conv.scala 25:31]
  assign conv_unit_1_io_bias2 = io_bias_data_3; // @[Conv.scala 26:31]
  assign conv_unit_1_io_bias_valid = io_bias_valid; // @[Conv.scala 27:36]
  assign conv_unit_2_clock = clock;
  assign conv_unit_2_io_ifm_win_33_0 = io_ifm_win_33_0; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_1 = io_ifm_win_33_1; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_2 = io_ifm_win_33_2; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_3 = io_ifm_win_33_3; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_4 = io_ifm_win_33_4; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_5 = io_ifm_win_33_5; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_6 = io_ifm_win_33_6; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_7 = io_ifm_win_33_7; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_8 = io_ifm_win_33_8; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_9 = io_ifm_win_33_9; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_10 = io_ifm_win_33_10; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_11 = io_ifm_win_33_11; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_12 = io_ifm_win_33_12; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_13 = io_ifm_win_33_13; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_14 = io_ifm_win_33_14; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_15 = io_ifm_win_33_15; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_16 = io_ifm_win_33_16; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_17 = io_ifm_win_33_17; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_18 = io_ifm_win_33_18; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_19 = io_ifm_win_33_19; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_20 = io_ifm_win_33_20; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_21 = io_ifm_win_33_21; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_22 = io_ifm_win_33_22; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_23 = io_ifm_win_33_23; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_24 = io_ifm_win_33_24; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_25 = io_ifm_win_33_25; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_26 = io_ifm_win_33_26; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_27 = io_ifm_win_33_27; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_28 = io_ifm_win_33_28; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_29 = io_ifm_win_33_29; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_30 = io_ifm_win_33_30; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_31 = io_ifm_win_33_31; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_32 = io_ifm_win_33_32; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_33 = io_ifm_win_33_33; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_34 = io_ifm_win_33_34; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_35 = io_ifm_win_33_35; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_36 = io_ifm_win_33_36; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_37 = io_ifm_win_33_37; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_38 = io_ifm_win_33_38; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_39 = io_ifm_win_33_39; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_40 = io_ifm_win_33_40; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_41 = io_ifm_win_33_41; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_42 = io_ifm_win_33_42; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_43 = io_ifm_win_33_43; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_44 = io_ifm_win_33_44; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_45 = io_ifm_win_33_45; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_46 = io_ifm_win_33_46; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_47 = io_ifm_win_33_47; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_48 = io_ifm_win_33_48; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_49 = io_ifm_win_33_49; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_50 = io_ifm_win_33_50; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_51 = io_ifm_win_33_51; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_52 = io_ifm_win_33_52; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_53 = io_ifm_win_33_53; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_54 = io_ifm_win_33_54; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_55 = io_ifm_win_33_55; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_56 = io_ifm_win_33_56; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_57 = io_ifm_win_33_57; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_58 = io_ifm_win_33_58; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_59 = io_ifm_win_33_59; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_60 = io_ifm_win_33_60; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_61 = io_ifm_win_33_61; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_62 = io_ifm_win_33_62; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_63 = io_ifm_win_33_63; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_64 = io_ifm_win_33_64; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_65 = io_ifm_win_33_65; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_66 = io_ifm_win_33_66; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_67 = io_ifm_win_33_67; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_68 = io_ifm_win_33_68; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_69 = io_ifm_win_33_69; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_70 = io_ifm_win_33_70; // @[Conv.scala 20:36]
  assign conv_unit_2_io_ifm_win_33_71 = io_ifm_win_33_71; // @[Conv.scala 20:36]
  assign conv_unit_2_io_weight_win_33_ch1_0 = io_weight_win_33_288; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_1 = io_weight_win_33_289; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_2 = io_weight_win_33_290; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_3 = io_weight_win_33_291; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_4 = io_weight_win_33_292; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_5 = io_weight_win_33_293; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_6 = io_weight_win_33_294; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_7 = io_weight_win_33_295; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_8 = io_weight_win_33_296; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_9 = io_weight_win_33_297; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_10 = io_weight_win_33_298; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_11 = io_weight_win_33_299; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_12 = io_weight_win_33_300; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_13 = io_weight_win_33_301; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_14 = io_weight_win_33_302; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_15 = io_weight_win_33_303; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_16 = io_weight_win_33_304; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_17 = io_weight_win_33_305; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_18 = io_weight_win_33_306; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_19 = io_weight_win_33_307; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_20 = io_weight_win_33_308; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_21 = io_weight_win_33_309; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_22 = io_weight_win_33_310; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_23 = io_weight_win_33_311; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_24 = io_weight_win_33_312; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_25 = io_weight_win_33_313; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_26 = io_weight_win_33_314; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_27 = io_weight_win_33_315; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_28 = io_weight_win_33_316; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_29 = io_weight_win_33_317; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_30 = io_weight_win_33_318; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_31 = io_weight_win_33_319; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_32 = io_weight_win_33_320; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_33 = io_weight_win_33_321; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_34 = io_weight_win_33_322; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_35 = io_weight_win_33_323; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_36 = io_weight_win_33_324; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_37 = io_weight_win_33_325; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_38 = io_weight_win_33_326; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_39 = io_weight_win_33_327; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_40 = io_weight_win_33_328; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_41 = io_weight_win_33_329; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_42 = io_weight_win_33_330; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_43 = io_weight_win_33_331; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_44 = io_weight_win_33_332; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_45 = io_weight_win_33_333; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_46 = io_weight_win_33_334; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_47 = io_weight_win_33_335; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_48 = io_weight_win_33_336; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_49 = io_weight_win_33_337; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_50 = io_weight_win_33_338; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_51 = io_weight_win_33_339; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_52 = io_weight_win_33_340; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_53 = io_weight_win_33_341; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_54 = io_weight_win_33_342; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_55 = io_weight_win_33_343; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_56 = io_weight_win_33_344; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_57 = io_weight_win_33_345; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_58 = io_weight_win_33_346; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_59 = io_weight_win_33_347; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_60 = io_weight_win_33_348; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_61 = io_weight_win_33_349; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_62 = io_weight_win_33_350; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_63 = io_weight_win_33_351; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_64 = io_weight_win_33_352; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_65 = io_weight_win_33_353; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_66 = io_weight_win_33_354; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_67 = io_weight_win_33_355; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_68 = io_weight_win_33_356; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_69 = io_weight_win_33_357; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_70 = io_weight_win_33_358; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch1_71 = io_weight_win_33_359; // @[Conv.scala 22:50]
  assign conv_unit_2_io_weight_win_33_ch2_0 = io_weight_win_33_360; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_1 = io_weight_win_33_361; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_2 = io_weight_win_33_362; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_3 = io_weight_win_33_363; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_4 = io_weight_win_33_364; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_5 = io_weight_win_33_365; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_6 = io_weight_win_33_366; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_7 = io_weight_win_33_367; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_8 = io_weight_win_33_368; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_9 = io_weight_win_33_369; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_10 = io_weight_win_33_370; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_11 = io_weight_win_33_371; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_12 = io_weight_win_33_372; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_13 = io_weight_win_33_373; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_14 = io_weight_win_33_374; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_15 = io_weight_win_33_375; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_16 = io_weight_win_33_376; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_17 = io_weight_win_33_377; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_18 = io_weight_win_33_378; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_19 = io_weight_win_33_379; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_20 = io_weight_win_33_380; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_21 = io_weight_win_33_381; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_22 = io_weight_win_33_382; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_23 = io_weight_win_33_383; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_24 = io_weight_win_33_384; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_25 = io_weight_win_33_385; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_26 = io_weight_win_33_386; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_27 = io_weight_win_33_387; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_28 = io_weight_win_33_388; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_29 = io_weight_win_33_389; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_30 = io_weight_win_33_390; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_31 = io_weight_win_33_391; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_32 = io_weight_win_33_392; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_33 = io_weight_win_33_393; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_34 = io_weight_win_33_394; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_35 = io_weight_win_33_395; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_36 = io_weight_win_33_396; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_37 = io_weight_win_33_397; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_38 = io_weight_win_33_398; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_39 = io_weight_win_33_399; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_40 = io_weight_win_33_400; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_41 = io_weight_win_33_401; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_42 = io_weight_win_33_402; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_43 = io_weight_win_33_403; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_44 = io_weight_win_33_404; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_45 = io_weight_win_33_405; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_46 = io_weight_win_33_406; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_47 = io_weight_win_33_407; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_48 = io_weight_win_33_408; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_49 = io_weight_win_33_409; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_50 = io_weight_win_33_410; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_51 = io_weight_win_33_411; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_52 = io_weight_win_33_412; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_53 = io_weight_win_33_413; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_54 = io_weight_win_33_414; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_55 = io_weight_win_33_415; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_56 = io_weight_win_33_416; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_57 = io_weight_win_33_417; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_58 = io_weight_win_33_418; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_59 = io_weight_win_33_419; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_60 = io_weight_win_33_420; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_61 = io_weight_win_33_421; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_62 = io_weight_win_33_422; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_63 = io_weight_win_33_423; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_64 = io_weight_win_33_424; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_65 = io_weight_win_33_425; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_66 = io_weight_win_33_426; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_67 = io_weight_win_33_427; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_68 = io_weight_win_33_428; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_69 = io_weight_win_33_429; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_70 = io_weight_win_33_430; // @[Conv.scala 23:50]
  assign conv_unit_2_io_weight_win_33_ch2_71 = io_weight_win_33_431; // @[Conv.scala 23:50]
  assign conv_unit_2_io_bias1 = io_bias_data_4; // @[Conv.scala 25:31]
  assign conv_unit_2_io_bias2 = io_bias_data_5; // @[Conv.scala 26:31]
  assign conv_unit_2_io_bias_valid = io_bias_valid; // @[Conv.scala 27:36]
  assign conv_unit_3_clock = clock;
  assign conv_unit_3_io_ifm_win_33_0 = io_ifm_win_33_0; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_1 = io_ifm_win_33_1; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_2 = io_ifm_win_33_2; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_3 = io_ifm_win_33_3; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_4 = io_ifm_win_33_4; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_5 = io_ifm_win_33_5; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_6 = io_ifm_win_33_6; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_7 = io_ifm_win_33_7; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_8 = io_ifm_win_33_8; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_9 = io_ifm_win_33_9; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_10 = io_ifm_win_33_10; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_11 = io_ifm_win_33_11; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_12 = io_ifm_win_33_12; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_13 = io_ifm_win_33_13; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_14 = io_ifm_win_33_14; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_15 = io_ifm_win_33_15; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_16 = io_ifm_win_33_16; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_17 = io_ifm_win_33_17; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_18 = io_ifm_win_33_18; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_19 = io_ifm_win_33_19; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_20 = io_ifm_win_33_20; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_21 = io_ifm_win_33_21; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_22 = io_ifm_win_33_22; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_23 = io_ifm_win_33_23; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_24 = io_ifm_win_33_24; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_25 = io_ifm_win_33_25; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_26 = io_ifm_win_33_26; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_27 = io_ifm_win_33_27; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_28 = io_ifm_win_33_28; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_29 = io_ifm_win_33_29; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_30 = io_ifm_win_33_30; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_31 = io_ifm_win_33_31; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_32 = io_ifm_win_33_32; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_33 = io_ifm_win_33_33; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_34 = io_ifm_win_33_34; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_35 = io_ifm_win_33_35; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_36 = io_ifm_win_33_36; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_37 = io_ifm_win_33_37; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_38 = io_ifm_win_33_38; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_39 = io_ifm_win_33_39; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_40 = io_ifm_win_33_40; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_41 = io_ifm_win_33_41; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_42 = io_ifm_win_33_42; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_43 = io_ifm_win_33_43; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_44 = io_ifm_win_33_44; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_45 = io_ifm_win_33_45; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_46 = io_ifm_win_33_46; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_47 = io_ifm_win_33_47; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_48 = io_ifm_win_33_48; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_49 = io_ifm_win_33_49; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_50 = io_ifm_win_33_50; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_51 = io_ifm_win_33_51; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_52 = io_ifm_win_33_52; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_53 = io_ifm_win_33_53; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_54 = io_ifm_win_33_54; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_55 = io_ifm_win_33_55; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_56 = io_ifm_win_33_56; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_57 = io_ifm_win_33_57; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_58 = io_ifm_win_33_58; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_59 = io_ifm_win_33_59; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_60 = io_ifm_win_33_60; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_61 = io_ifm_win_33_61; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_62 = io_ifm_win_33_62; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_63 = io_ifm_win_33_63; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_64 = io_ifm_win_33_64; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_65 = io_ifm_win_33_65; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_66 = io_ifm_win_33_66; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_67 = io_ifm_win_33_67; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_68 = io_ifm_win_33_68; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_69 = io_ifm_win_33_69; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_70 = io_ifm_win_33_70; // @[Conv.scala 20:36]
  assign conv_unit_3_io_ifm_win_33_71 = io_ifm_win_33_71; // @[Conv.scala 20:36]
  assign conv_unit_3_io_weight_win_33_ch1_0 = io_weight_win_33_432; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_1 = io_weight_win_33_433; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_2 = io_weight_win_33_434; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_3 = io_weight_win_33_435; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_4 = io_weight_win_33_436; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_5 = io_weight_win_33_437; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_6 = io_weight_win_33_438; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_7 = io_weight_win_33_439; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_8 = io_weight_win_33_440; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_9 = io_weight_win_33_441; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_10 = io_weight_win_33_442; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_11 = io_weight_win_33_443; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_12 = io_weight_win_33_444; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_13 = io_weight_win_33_445; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_14 = io_weight_win_33_446; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_15 = io_weight_win_33_447; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_16 = io_weight_win_33_448; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_17 = io_weight_win_33_449; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_18 = io_weight_win_33_450; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_19 = io_weight_win_33_451; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_20 = io_weight_win_33_452; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_21 = io_weight_win_33_453; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_22 = io_weight_win_33_454; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_23 = io_weight_win_33_455; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_24 = io_weight_win_33_456; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_25 = io_weight_win_33_457; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_26 = io_weight_win_33_458; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_27 = io_weight_win_33_459; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_28 = io_weight_win_33_460; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_29 = io_weight_win_33_461; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_30 = io_weight_win_33_462; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_31 = io_weight_win_33_463; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_32 = io_weight_win_33_464; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_33 = io_weight_win_33_465; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_34 = io_weight_win_33_466; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_35 = io_weight_win_33_467; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_36 = io_weight_win_33_468; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_37 = io_weight_win_33_469; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_38 = io_weight_win_33_470; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_39 = io_weight_win_33_471; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_40 = io_weight_win_33_472; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_41 = io_weight_win_33_473; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_42 = io_weight_win_33_474; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_43 = io_weight_win_33_475; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_44 = io_weight_win_33_476; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_45 = io_weight_win_33_477; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_46 = io_weight_win_33_478; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_47 = io_weight_win_33_479; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_48 = io_weight_win_33_480; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_49 = io_weight_win_33_481; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_50 = io_weight_win_33_482; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_51 = io_weight_win_33_483; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_52 = io_weight_win_33_484; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_53 = io_weight_win_33_485; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_54 = io_weight_win_33_486; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_55 = io_weight_win_33_487; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_56 = io_weight_win_33_488; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_57 = io_weight_win_33_489; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_58 = io_weight_win_33_490; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_59 = io_weight_win_33_491; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_60 = io_weight_win_33_492; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_61 = io_weight_win_33_493; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_62 = io_weight_win_33_494; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_63 = io_weight_win_33_495; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_64 = io_weight_win_33_496; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_65 = io_weight_win_33_497; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_66 = io_weight_win_33_498; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_67 = io_weight_win_33_499; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_68 = io_weight_win_33_500; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_69 = io_weight_win_33_501; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_70 = io_weight_win_33_502; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch1_71 = io_weight_win_33_503; // @[Conv.scala 22:50]
  assign conv_unit_3_io_weight_win_33_ch2_0 = io_weight_win_33_504; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_1 = io_weight_win_33_505; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_2 = io_weight_win_33_506; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_3 = io_weight_win_33_507; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_4 = io_weight_win_33_508; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_5 = io_weight_win_33_509; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_6 = io_weight_win_33_510; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_7 = io_weight_win_33_511; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_8 = io_weight_win_33_512; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_9 = io_weight_win_33_513; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_10 = io_weight_win_33_514; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_11 = io_weight_win_33_515; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_12 = io_weight_win_33_516; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_13 = io_weight_win_33_517; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_14 = io_weight_win_33_518; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_15 = io_weight_win_33_519; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_16 = io_weight_win_33_520; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_17 = io_weight_win_33_521; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_18 = io_weight_win_33_522; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_19 = io_weight_win_33_523; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_20 = io_weight_win_33_524; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_21 = io_weight_win_33_525; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_22 = io_weight_win_33_526; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_23 = io_weight_win_33_527; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_24 = io_weight_win_33_528; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_25 = io_weight_win_33_529; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_26 = io_weight_win_33_530; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_27 = io_weight_win_33_531; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_28 = io_weight_win_33_532; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_29 = io_weight_win_33_533; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_30 = io_weight_win_33_534; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_31 = io_weight_win_33_535; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_32 = io_weight_win_33_536; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_33 = io_weight_win_33_537; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_34 = io_weight_win_33_538; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_35 = io_weight_win_33_539; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_36 = io_weight_win_33_540; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_37 = io_weight_win_33_541; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_38 = io_weight_win_33_542; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_39 = io_weight_win_33_543; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_40 = io_weight_win_33_544; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_41 = io_weight_win_33_545; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_42 = io_weight_win_33_546; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_43 = io_weight_win_33_547; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_44 = io_weight_win_33_548; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_45 = io_weight_win_33_549; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_46 = io_weight_win_33_550; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_47 = io_weight_win_33_551; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_48 = io_weight_win_33_552; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_49 = io_weight_win_33_553; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_50 = io_weight_win_33_554; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_51 = io_weight_win_33_555; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_52 = io_weight_win_33_556; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_53 = io_weight_win_33_557; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_54 = io_weight_win_33_558; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_55 = io_weight_win_33_559; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_56 = io_weight_win_33_560; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_57 = io_weight_win_33_561; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_58 = io_weight_win_33_562; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_59 = io_weight_win_33_563; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_60 = io_weight_win_33_564; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_61 = io_weight_win_33_565; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_62 = io_weight_win_33_566; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_63 = io_weight_win_33_567; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_64 = io_weight_win_33_568; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_65 = io_weight_win_33_569; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_66 = io_weight_win_33_570; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_67 = io_weight_win_33_571; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_68 = io_weight_win_33_572; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_69 = io_weight_win_33_573; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_70 = io_weight_win_33_574; // @[Conv.scala 23:50]
  assign conv_unit_3_io_weight_win_33_ch2_71 = io_weight_win_33_575; // @[Conv.scala 23:50]
  assign conv_unit_3_io_bias1 = io_bias_data_6; // @[Conv.scala 25:31]
  assign conv_unit_3_io_bias2 = io_bias_data_7; // @[Conv.scala 26:31]
  assign conv_unit_3_io_bias_valid = io_bias_valid; // @[Conv.scala 27:36]
endmodule
module TPRAM_WRAP_88(
  input         clock,
  input         io_wen,
  input         io_ren,
  input  [11:0] io_waddr,
  input  [11:0] io_raddr,
  input  [17:0] io_wdata,
  output [17:0] io_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  tpram_CLKA; // @[utils.scala 218:23]
  wire  tpram_CLKB; // @[utils.scala 218:23]
  wire  tpram_CENB; // @[utils.scala 218:23]
  wire  tpram_CENA; // @[utils.scala 218:23]
  wire [11:0] tpram_AB; // @[utils.scala 218:23]
  wire [11:0] tpram_AA; // @[utils.scala 218:23]
  wire [17:0] tpram_DB; // @[utils.scala 218:23]
  wire [17:0] tpram_QA; // @[utils.scala 218:23]
  reg  rd_en; // @[utils.scala 219:46]
  reg [17:0] rdata_reg; // @[Reg.scala 19:16]
  TPRAM #(.DATA_WIDTH(18), .DEPTH(4096), .RAM_STYLE_VAL("block")) tpram ( // @[utils.scala 218:23]
    .CLKA(tpram_CLKA),
    .CLKB(tpram_CLKB),
    .CENB(tpram_CENB),
    .CENA(tpram_CENA),
    .AB(tpram_AB),
    .AA(tpram_AA),
    .DB(tpram_DB),
    .QA(tpram_QA)
  );
  assign io_rdata = ~rd_en ? rdata_reg : tpram_QA; // @[utils.scala 230:12]
  assign tpram_CLKA = clock; // @[utils.scala 222:19]
  assign tpram_CLKB = clock; // @[utils.scala 223:19]
  assign tpram_CENB = ~io_wen; // @[utils.scala 224:22]
  assign tpram_CENA = ~io_ren; // @[utils.scala 225:22]
  assign tpram_AB = io_waddr; // @[utils.scala 226:17]
  assign tpram_AA = io_raddr; // @[utils.scala 227:17]
  assign tpram_DB = io_wdata; // @[utils.scala 228:17]
  always @(posedge clock) begin
    rd_en <= io_ren; // @[utils.scala 219:46]
    if (rd_en) begin // @[Reg.scala 20:18]
      rdata_reg <= tpram_QA; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rd_en = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rdata_reg = _RAND_1[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cal_acc_unit(
  input         clock,
  input         reset,
  input  [17:0] io_a,
  input  [17:0] io_b,
  input         io_a_zero,
  input         io_b_zero,
  output [17:0] io_c
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] c_t; // @[utils.scala 850:22]
  wire [17:0] a_z = io_a_zero ? $signed(18'sh0) : $signed(io_a); // @[utils.scala 851:15]
  wire [17:0] b_z = io_b_zero ? $signed(18'sh0) : $signed(io_b); // @[utils.scala 852:15]
  wire [17:0] _c_t_T_2 = $signed(a_z) + $signed(b_z); // @[utils.scala 853:16]
  assign io_c = c_t; // @[utils.scala 854:10]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 850:22]
      c_t <= 18'sh0; // @[utils.scala 850:22]
    end else begin
      c_t <= _c_t_T_2; // @[utils.scala 853:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  c_t = _RAND_0[17:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module acc_mem_unit(
  input         clock,
  input         reset,
  input         io_prev_data_zero,
  input         io_curr_data_zero,
  input         io_read_en,
  input         io_write_en,
  input  [11:0] io_read_addr,
  input  [11:0] io_write_addr,
  input  [17:0] io_curr_data,
  output [17:0] io_acc_result
);
  wire  TPRAM_WRAP_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_wen; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_ren; // @[utils.scala 237:100]
  wire [11:0] TPRAM_WRAP_io_waddr; // @[utils.scala 237:100]
  wire [11:0] TPRAM_WRAP_io_raddr; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_io_wdata; // @[utils.scala 237:100]
  wire [17:0] TPRAM_WRAP_io_rdata; // @[utils.scala 237:100]
  wire  acc_clock; // @[acc_mem.scala 55:21]
  wire  acc_reset; // @[acc_mem.scala 55:21]
  wire [17:0] acc_io_a; // @[acc_mem.scala 55:21]
  wire [17:0] acc_io_b; // @[acc_mem.scala 55:21]
  wire  acc_io_a_zero; // @[acc_mem.scala 55:21]
  wire  acc_io_b_zero; // @[acc_mem.scala 55:21]
  wire [17:0] acc_io_c; // @[acc_mem.scala 55:21]
  TPRAM_WRAP_88 TPRAM_WRAP ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_clock),
    .io_wen(TPRAM_WRAP_io_wen),
    .io_ren(TPRAM_WRAP_io_ren),
    .io_waddr(TPRAM_WRAP_io_waddr),
    .io_raddr(TPRAM_WRAP_io_raddr),
    .io_wdata(TPRAM_WRAP_io_wdata),
    .io_rdata(TPRAM_WRAP_io_rdata)
  );
  cal_acc_unit acc ( // @[acc_mem.scala 55:21]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_a(acc_io_a),
    .io_b(acc_io_b),
    .io_a_zero(acc_io_a_zero),
    .io_b_zero(acc_io_b_zero),
    .io_c(acc_io_c)
  );
  assign io_acc_result = acc_io_c; // @[acc_mem.scala 60:27]
  assign TPRAM_WRAP_clock = clock;
  assign TPRAM_WRAP_io_wen = io_write_en; // @[acc_mem.scala 48:13]
  assign TPRAM_WRAP_io_ren = io_read_en; // @[acc_mem.scala 49:13]
  assign TPRAM_WRAP_io_waddr = io_write_addr; // @[acc_mem.scala 50:15]
  assign TPRAM_WRAP_io_raddr = io_read_addr; // @[acc_mem.scala 51:15]
  assign TPRAM_WRAP_io_wdata = acc_io_c; // @[acc_mem.scala 60:27]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_a = TPRAM_WRAP_io_rdata; // @[acc_mem.scala 58:27]
  assign acc_io_b = io_curr_data; // @[acc_mem.scala 59:30]
  assign acc_io_a_zero = io_prev_data_zero; // @[acc_mem.scala 56:19]
  assign acc_io_b_zero = io_curr_data_zero; // @[acc_mem.scala 57:19]
endmodule
module acc(
  input         clock,
  input         reset,
  input         io_prev_data_zero,
  input         io_curr_data_zero,
  input         io_read_en,
  input         io_write_en,
  input  [11:0] io_read_addr,
  input  [11:0] io_write_addr,
  input  [17:0] io_curr_data_0,
  input  [17:0] io_curr_data_1,
  input  [17:0] io_curr_data_2,
  input  [17:0] io_curr_data_3,
  input  [17:0] io_curr_data_4,
  input  [17:0] io_curr_data_5,
  input  [17:0] io_curr_data_6,
  input  [17:0] io_curr_data_7,
  output [17:0] io_acc_result_0,
  output [17:0] io_acc_result_1,
  output [17:0] io_acc_result_2,
  output [17:0] io_acc_result_3,
  output [17:0] io_acc_result_4,
  output [17:0] io_acc_result_5,
  output [17:0] io_acc_result_6,
  output [17:0] io_acc_result_7
);
  wire  acc_unit_0_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_0_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_0_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_0_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_0_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_0_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_0_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_0_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_0_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_0_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_1_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_1_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_1_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_1_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_1_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_2_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_2_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_2_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_2_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_2_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_3_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_3_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_3_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_3_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_3_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_4_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_4_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_4_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_4_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_4_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_5_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_5_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_5_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_5_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_5_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_6_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_6_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_6_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_6_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_6_io_acc_result; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_clock; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_reset; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_io_prev_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_io_curr_data_zero; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_io_read_en; // @[acc_mem.scala 19:42]
  wire  acc_unit_7_io_write_en; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_7_io_read_addr; // @[acc_mem.scala 19:42]
  wire [11:0] acc_unit_7_io_write_addr; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_7_io_curr_data; // @[acc_mem.scala 19:42]
  wire [17:0] acc_unit_7_io_acc_result; // @[acc_mem.scala 19:42]
  acc_mem_unit acc_unit_0 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_0_clock),
    .reset(acc_unit_0_reset),
    .io_prev_data_zero(acc_unit_0_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_0_io_curr_data_zero),
    .io_read_en(acc_unit_0_io_read_en),
    .io_write_en(acc_unit_0_io_write_en),
    .io_read_addr(acc_unit_0_io_read_addr),
    .io_write_addr(acc_unit_0_io_write_addr),
    .io_curr_data(acc_unit_0_io_curr_data),
    .io_acc_result(acc_unit_0_io_acc_result)
  );
  acc_mem_unit acc_unit_1 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_1_clock),
    .reset(acc_unit_1_reset),
    .io_prev_data_zero(acc_unit_1_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_1_io_curr_data_zero),
    .io_read_en(acc_unit_1_io_read_en),
    .io_write_en(acc_unit_1_io_write_en),
    .io_read_addr(acc_unit_1_io_read_addr),
    .io_write_addr(acc_unit_1_io_write_addr),
    .io_curr_data(acc_unit_1_io_curr_data),
    .io_acc_result(acc_unit_1_io_acc_result)
  );
  acc_mem_unit acc_unit_2 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_2_clock),
    .reset(acc_unit_2_reset),
    .io_prev_data_zero(acc_unit_2_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_2_io_curr_data_zero),
    .io_read_en(acc_unit_2_io_read_en),
    .io_write_en(acc_unit_2_io_write_en),
    .io_read_addr(acc_unit_2_io_read_addr),
    .io_write_addr(acc_unit_2_io_write_addr),
    .io_curr_data(acc_unit_2_io_curr_data),
    .io_acc_result(acc_unit_2_io_acc_result)
  );
  acc_mem_unit acc_unit_3 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_3_clock),
    .reset(acc_unit_3_reset),
    .io_prev_data_zero(acc_unit_3_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_3_io_curr_data_zero),
    .io_read_en(acc_unit_3_io_read_en),
    .io_write_en(acc_unit_3_io_write_en),
    .io_read_addr(acc_unit_3_io_read_addr),
    .io_write_addr(acc_unit_3_io_write_addr),
    .io_curr_data(acc_unit_3_io_curr_data),
    .io_acc_result(acc_unit_3_io_acc_result)
  );
  acc_mem_unit acc_unit_4 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_4_clock),
    .reset(acc_unit_4_reset),
    .io_prev_data_zero(acc_unit_4_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_4_io_curr_data_zero),
    .io_read_en(acc_unit_4_io_read_en),
    .io_write_en(acc_unit_4_io_write_en),
    .io_read_addr(acc_unit_4_io_read_addr),
    .io_write_addr(acc_unit_4_io_write_addr),
    .io_curr_data(acc_unit_4_io_curr_data),
    .io_acc_result(acc_unit_4_io_acc_result)
  );
  acc_mem_unit acc_unit_5 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_5_clock),
    .reset(acc_unit_5_reset),
    .io_prev_data_zero(acc_unit_5_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_5_io_curr_data_zero),
    .io_read_en(acc_unit_5_io_read_en),
    .io_write_en(acc_unit_5_io_write_en),
    .io_read_addr(acc_unit_5_io_read_addr),
    .io_write_addr(acc_unit_5_io_write_addr),
    .io_curr_data(acc_unit_5_io_curr_data),
    .io_acc_result(acc_unit_5_io_acc_result)
  );
  acc_mem_unit acc_unit_6 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_6_clock),
    .reset(acc_unit_6_reset),
    .io_prev_data_zero(acc_unit_6_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_6_io_curr_data_zero),
    .io_read_en(acc_unit_6_io_read_en),
    .io_write_en(acc_unit_6_io_write_en),
    .io_read_addr(acc_unit_6_io_read_addr),
    .io_write_addr(acc_unit_6_io_write_addr),
    .io_curr_data(acc_unit_6_io_curr_data),
    .io_acc_result(acc_unit_6_io_acc_result)
  );
  acc_mem_unit acc_unit_7 ( // @[acc_mem.scala 19:42]
    .clock(acc_unit_7_clock),
    .reset(acc_unit_7_reset),
    .io_prev_data_zero(acc_unit_7_io_prev_data_zero),
    .io_curr_data_zero(acc_unit_7_io_curr_data_zero),
    .io_read_en(acc_unit_7_io_read_en),
    .io_write_en(acc_unit_7_io_write_en),
    .io_read_addr(acc_unit_7_io_read_addr),
    .io_write_addr(acc_unit_7_io_write_addr),
    .io_curr_data(acc_unit_7_io_curr_data),
    .io_acc_result(acc_unit_7_io_acc_result)
  );
  assign io_acc_result_0 = acc_unit_0_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_1 = acc_unit_1_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_2 = acc_unit_2_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_3 = acc_unit_3_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_4 = acc_unit_4_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_5 = acc_unit_5_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_6 = acc_unit_6_io_acc_result; // @[acc_mem.scala 28:26]
  assign io_acc_result_7 = acc_unit_7_io_acc_result; // @[acc_mem.scala 28:26]
  assign acc_unit_0_clock = clock;
  assign acc_unit_0_reset = reset;
  assign acc_unit_0_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_0_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_0_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_0_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_0_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_0_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_0_io_curr_data = io_curr_data_0; // @[acc_mem.scala 27:34]
  assign acc_unit_1_clock = clock;
  assign acc_unit_1_reset = reset;
  assign acc_unit_1_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_1_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_1_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_1_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_1_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_1_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_1_io_curr_data = io_curr_data_1; // @[acc_mem.scala 27:34]
  assign acc_unit_2_clock = clock;
  assign acc_unit_2_reset = reset;
  assign acc_unit_2_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_2_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_2_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_2_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_2_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_2_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_2_io_curr_data = io_curr_data_2; // @[acc_mem.scala 27:34]
  assign acc_unit_3_clock = clock;
  assign acc_unit_3_reset = reset;
  assign acc_unit_3_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_3_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_3_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_3_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_3_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_3_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_3_io_curr_data = io_curr_data_3; // @[acc_mem.scala 27:34]
  assign acc_unit_4_clock = clock;
  assign acc_unit_4_reset = reset;
  assign acc_unit_4_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_4_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_4_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_4_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_4_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_4_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_4_io_curr_data = io_curr_data_4; // @[acc_mem.scala 27:34]
  assign acc_unit_5_clock = clock;
  assign acc_unit_5_reset = reset;
  assign acc_unit_5_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_5_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_5_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_5_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_5_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_5_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_5_io_curr_data = io_curr_data_5; // @[acc_mem.scala 27:34]
  assign acc_unit_6_clock = clock;
  assign acc_unit_6_reset = reset;
  assign acc_unit_6_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_6_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_6_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_6_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_6_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_6_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_6_io_curr_data = io_curr_data_6; // @[acc_mem.scala 27:34]
  assign acc_unit_7_clock = clock;
  assign acc_unit_7_reset = reset;
  assign acc_unit_7_io_prev_data_zero = io_prev_data_zero; // @[acc_mem.scala 21:39]
  assign acc_unit_7_io_curr_data_zero = io_curr_data_zero; // @[acc_mem.scala 22:39]
  assign acc_unit_7_io_read_en = io_read_en; // @[acc_mem.scala 23:32]
  assign acc_unit_7_io_write_en = io_write_en; // @[acc_mem.scala 24:33]
  assign acc_unit_7_io_read_addr = io_read_addr; // @[acc_mem.scala 25:34]
  assign acc_unit_7_io_write_addr = io_write_addr; // @[acc_mem.scala 26:35]
  assign acc_unit_7_io_curr_data = io_curr_data_7; // @[acc_mem.scala 27:34]
endmodule
module sat_int18_16(
  input         clock,
  input  [17:0] io_data_in,
  output [15:0] io_data_out
);
  wire  sat_clk; // @[utils.scala 756:21]
  wire [17:0] sat_data_in; // @[utils.scala 756:21]
  wire [15:0] sat_data_out; // @[utils.scala 756:21]
  cal_sat_int18_int16 sat ( // @[utils.scala 756:21]
    .clk(sat_clk),
    .data_in(sat_data_in),
    .data_out(sat_data_out)
  );
  assign io_data_out = sat_data_out; // @[utils.scala 759:17]
  assign sat_clk = clock; // @[utils.scala 757:16]
  assign sat_data_in = io_data_in; // @[utils.scala 758:20]
endmodule
module scale_mul(
  input         clock,
  input  [15:0] io_v,
  input  [15:0] io_scale,
  output [31:0] io_dout
);
  wire  m_clk; // @[utils.scala 798:19]
  wire [15:0] m_val_in; // @[utils.scala 798:19]
  wire [15:0] m_scale; // @[utils.scala 798:19]
  wire [31:0] m_dout; // @[utils.scala 798:19]
  cal_scale_mul m ( // @[utils.scala 798:19]
    .clk(m_clk),
    .val_in(m_val_in),
    .scale(m_scale),
    .dout(m_dout)
  );
  assign io_dout = m_dout; // @[utils.scala 802:13]
  assign m_clk = clock; // @[utils.scala 799:14]
  assign m_val_in = io_v; // @[utils.scala 800:17]
  assign m_scale = io_scale; // @[utils.scala 801:16]
endmodule
module scale_shift(
  input         clock,
  input  [31:0] io_din,
  input  [3:0]  io_shift,
  output [15:0] io_dout
);
  wire  m_clk; // @[utils.scala 821:19]
  wire [31:0] m_din; // @[utils.scala 821:19]
  wire [3:0] m_shift; // @[utils.scala 821:19]
  wire [15:0] m_dout; // @[utils.scala 821:19]
  cal_scale_shift m ( // @[utils.scala 821:19]
    .clk(m_clk),
    .din(m_din),
    .shift(m_shift),
    .dout(m_dout)
  );
  assign io_dout = m_dout; // @[utils.scala 825:13]
  assign m_clk = clock; // @[utils.scala 822:14]
  assign m_din = io_din; // @[utils.scala 823:14]
  assign m_shift = io_shift; // @[utils.scala 824:16]
endmodule
module scale(
  input         clock,
  input  [15:0] io_v,
  input  [15:0] io_scale,
  input  [3:0]  io_shift,
  output [15:0] io_dout
);
  wire  mul_clock; // @[quant.scala 62:21]
  wire [15:0] mul_io_v; // @[quant.scala 62:21]
  wire [15:0] mul_io_scale; // @[quant.scala 62:21]
  wire [31:0] mul_io_dout; // @[quant.scala 62:21]
  wire  shift_clock; // @[quant.scala 66:23]
  wire [31:0] shift_io_din; // @[quant.scala 66:23]
  wire [3:0] shift_io_shift; // @[quant.scala 66:23]
  wire [15:0] shift_io_dout; // @[quant.scala 66:23]
  scale_mul mul ( // @[quant.scala 62:21]
    .clock(mul_clock),
    .io_v(mul_io_v),
    .io_scale(mul_io_scale),
    .io_dout(mul_io_dout)
  );
  scale_shift shift ( // @[quant.scala 66:23]
    .clock(shift_clock),
    .io_din(shift_io_din),
    .io_shift(shift_io_shift),
    .io_dout(shift_io_dout)
  );
  assign io_dout = shift_io_dout; // @[quant.scala 69:13]
  assign mul_clock = clock;
  assign mul_io_v = io_v; // @[quant.scala 63:14]
  assign mul_io_scale = io_scale; // @[quant.scala 64:18]
  assign shift_clock = clock;
  assign shift_io_din = mul_io_dout; // @[quant.scala 61:20 65:10]
  assign shift_io_shift = io_shift; // @[quant.scala 68:20]
endmodule
module sat_int16_8(
  input         clock,
  input  [15:0] io_data_in,
  output [7:0]  io_data_out
);
  wire  sat_clk; // @[utils.scala 776:21]
  wire [15:0] sat_data_in; // @[utils.scala 776:21]
  wire [7:0] sat_data_out; // @[utils.scala 776:21]
  cal_sat_int16_int8 sat ( // @[utils.scala 776:21]
    .clk(sat_clk),
    .data_in(sat_data_in),
    .data_out(sat_data_out)
  );
  assign io_data_out = sat_data_out; // @[utils.scala 779:17]
  assign sat_clk = clock; // @[utils.scala 777:16]
  assign sat_data_in = io_data_in; // @[utils.scala 778:20]
endmodule
module quant_unit(
  input         clock,
  input  [17:0] io_acc_result,
  input  [15:0] io_scale,
  input  [3:0]  io_shift,
  input  [7:0]  io_zero_point,
  output [7:0]  io_quant_result
);
  wire  sat_18_16_clock; // @[quant.scala 36:27]
  wire [17:0] sat_18_16_io_data_in; // @[quant.scala 36:27]
  wire [15:0] sat_18_16_io_data_out; // @[quant.scala 36:27]
  wire  scale_clock; // @[quant.scala 40:23]
  wire [15:0] scale_io_v; // @[quant.scala 40:23]
  wire [15:0] scale_io_scale; // @[quant.scala 40:23]
  wire [3:0] scale_io_shift; // @[quant.scala 40:23]
  wire [15:0] scale_io_dout; // @[quant.scala 40:23]
  wire  sat_16_8_clock; // @[quant.scala 46:26]
  wire [15:0] sat_16_8_io_data_in; // @[quant.scala 46:26]
  wire [7:0] sat_16_8_io_data_out; // @[quant.scala 46:26]
  wire [7:0] _after_sat8_T = sat_16_8_io_data_out; // @[quant.scala 48:40]
  wire [7:0] _temp_T = io_zero_point; // @[quant.scala 50:43]
  wire [15:0] after_sat8 = {{8{_after_sat8_T[7]}},_after_sat8_T}; // @[quant.scala 34:26 48:16]
  wire [15:0] _GEN_0 = {{8{_temp_T[7]}},_temp_T}; // @[quant.scala 50:27]
  wire [15:0] _io_quant_result_T = $signed(after_sat8) + $signed(_GEN_0); // @[quant.scala 51:29]
  sat_int18_16 sat_18_16 ( // @[quant.scala 36:27]
    .clock(sat_18_16_clock),
    .io_data_in(sat_18_16_io_data_in),
    .io_data_out(sat_18_16_io_data_out)
  );
  scale scale ( // @[quant.scala 40:23]
    .clock(scale_clock),
    .io_v(scale_io_v),
    .io_scale(scale_io_scale),
    .io_shift(scale_io_shift),
    .io_dout(scale_io_dout)
  );
  sat_int16_8 sat_16_8 ( // @[quant.scala 46:26]
    .clock(sat_16_8_clock),
    .io_data_in(sat_16_8_io_data_in),
    .io_data_out(sat_16_8_io_data_out)
  );
  assign io_quant_result = _io_quant_result_T[7:0]; // @[quant.scala 51:21]
  assign sat_18_16_clock = clock;
  assign sat_18_16_io_data_in = io_acc_result; // @[quant.scala 37:26]
  assign scale_clock = clock;
  assign scale_io_v = sat_18_16_io_data_out; // @[quant.scala 41:35]
  assign scale_io_scale = io_scale; // @[quant.scala 42:32]
  assign scale_io_shift = io_shift; // @[quant.scala 43:20]
  assign sat_16_8_clock = clock;
  assign sat_16_8_io_data_in = scale_io_dout; // @[quant.scala 44:34]
endmodule
module quant(
  input         clock,
  input  [17:0] io_acc_result_0,
  input  [17:0] io_acc_result_1,
  input  [17:0] io_acc_result_2,
  input  [17:0] io_acc_result_3,
  input  [17:0] io_acc_result_4,
  input  [17:0] io_acc_result_5,
  input  [17:0] io_acc_result_6,
  input  [17:0] io_acc_result_7,
  input  [15:0] io_scale,
  input  [3:0]  io_shift,
  input  [7:0]  io_zero_point,
  output [7:0]  io_quant_result_0,
  output [7:0]  io_quant_result_1,
  output [7:0]  io_quant_result_2,
  output [7:0]  io_quant_result_3,
  output [7:0]  io_quant_result_4,
  output [7:0]  io_quant_result_5,
  output [7:0]  io_quant_result_6,
  output [7:0]  io_quant_result_7
);
  wire  quant_unit_0_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_0_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_0_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_0_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_0_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_0_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_1_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_1_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_1_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_1_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_1_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_1_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_2_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_2_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_2_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_2_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_2_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_2_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_3_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_3_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_3_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_3_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_3_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_3_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_4_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_4_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_4_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_4_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_4_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_4_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_5_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_5_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_5_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_5_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_5_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_5_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_6_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_6_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_6_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_6_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_6_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_6_io_quant_result; // @[quant.scala 14:56]
  wire  quant_unit_7_clock; // @[quant.scala 14:56]
  wire [17:0] quant_unit_7_io_acc_result; // @[quant.scala 14:56]
  wire [15:0] quant_unit_7_io_scale; // @[quant.scala 14:56]
  wire [3:0] quant_unit_7_io_shift; // @[quant.scala 14:56]
  wire [7:0] quant_unit_7_io_zero_point; // @[quant.scala 14:56]
  wire [7:0] quant_unit_7_io_quant_result; // @[quant.scala 14:56]
  quant_unit quant_unit_0 ( // @[quant.scala 14:56]
    .clock(quant_unit_0_clock),
    .io_acc_result(quant_unit_0_io_acc_result),
    .io_scale(quant_unit_0_io_scale),
    .io_shift(quant_unit_0_io_shift),
    .io_zero_point(quant_unit_0_io_zero_point),
    .io_quant_result(quant_unit_0_io_quant_result)
  );
  quant_unit quant_unit_1 ( // @[quant.scala 14:56]
    .clock(quant_unit_1_clock),
    .io_acc_result(quant_unit_1_io_acc_result),
    .io_scale(quant_unit_1_io_scale),
    .io_shift(quant_unit_1_io_shift),
    .io_zero_point(quant_unit_1_io_zero_point),
    .io_quant_result(quant_unit_1_io_quant_result)
  );
  quant_unit quant_unit_2 ( // @[quant.scala 14:56]
    .clock(quant_unit_2_clock),
    .io_acc_result(quant_unit_2_io_acc_result),
    .io_scale(quant_unit_2_io_scale),
    .io_shift(quant_unit_2_io_shift),
    .io_zero_point(quant_unit_2_io_zero_point),
    .io_quant_result(quant_unit_2_io_quant_result)
  );
  quant_unit quant_unit_3 ( // @[quant.scala 14:56]
    .clock(quant_unit_3_clock),
    .io_acc_result(quant_unit_3_io_acc_result),
    .io_scale(quant_unit_3_io_scale),
    .io_shift(quant_unit_3_io_shift),
    .io_zero_point(quant_unit_3_io_zero_point),
    .io_quant_result(quant_unit_3_io_quant_result)
  );
  quant_unit quant_unit_4 ( // @[quant.scala 14:56]
    .clock(quant_unit_4_clock),
    .io_acc_result(quant_unit_4_io_acc_result),
    .io_scale(quant_unit_4_io_scale),
    .io_shift(quant_unit_4_io_shift),
    .io_zero_point(quant_unit_4_io_zero_point),
    .io_quant_result(quant_unit_4_io_quant_result)
  );
  quant_unit quant_unit_5 ( // @[quant.scala 14:56]
    .clock(quant_unit_5_clock),
    .io_acc_result(quant_unit_5_io_acc_result),
    .io_scale(quant_unit_5_io_scale),
    .io_shift(quant_unit_5_io_shift),
    .io_zero_point(quant_unit_5_io_zero_point),
    .io_quant_result(quant_unit_5_io_quant_result)
  );
  quant_unit quant_unit_6 ( // @[quant.scala 14:56]
    .clock(quant_unit_6_clock),
    .io_acc_result(quant_unit_6_io_acc_result),
    .io_scale(quant_unit_6_io_scale),
    .io_shift(quant_unit_6_io_shift),
    .io_zero_point(quant_unit_6_io_zero_point),
    .io_quant_result(quant_unit_6_io_quant_result)
  );
  quant_unit quant_unit_7 ( // @[quant.scala 14:56]
    .clock(quant_unit_7_clock),
    .io_acc_result(quant_unit_7_io_acc_result),
    .io_scale(quant_unit_7_io_scale),
    .io_shift(quant_unit_7_io_shift),
    .io_zero_point(quant_unit_7_io_zero_point),
    .io_quant_result(quant_unit_7_io_quant_result)
  );
  assign io_quant_result_0 = quant_unit_0_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_1 = quant_unit_1_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_2 = quant_unit_2_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_3 = quant_unit_3_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_4 = quant_unit_4_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_5 = quant_unit_5_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_6 = quant_unit_6_io_quant_result; // @[quant.scala 20:28]
  assign io_quant_result_7 = quant_unit_7_io_quant_result; // @[quant.scala 20:28]
  assign quant_unit_0_clock = clock;
  assign quant_unit_0_io_acc_result = io_acc_result_0; // @[quant.scala 16:37]
  assign quant_unit_0_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_0_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_0_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_1_clock = clock;
  assign quant_unit_1_io_acc_result = io_acc_result_1; // @[quant.scala 16:37]
  assign quant_unit_1_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_1_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_1_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_2_clock = clock;
  assign quant_unit_2_io_acc_result = io_acc_result_2; // @[quant.scala 16:37]
  assign quant_unit_2_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_2_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_2_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_3_clock = clock;
  assign quant_unit_3_io_acc_result = io_acc_result_3; // @[quant.scala 16:37]
  assign quant_unit_3_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_3_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_3_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_4_clock = clock;
  assign quant_unit_4_io_acc_result = io_acc_result_4; // @[quant.scala 16:37]
  assign quant_unit_4_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_4_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_4_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_5_clock = clock;
  assign quant_unit_5_io_acc_result = io_acc_result_5; // @[quant.scala 16:37]
  assign quant_unit_5_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_5_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_5_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_6_clock = clock;
  assign quant_unit_6_io_acc_result = io_acc_result_6; // @[quant.scala 16:37]
  assign quant_unit_6_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_6_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_6_io_zero_point = io_zero_point; // @[quant.scala 19:37]
  assign quant_unit_7_clock = clock;
  assign quant_unit_7_io_acc_result = io_acc_result_7; // @[quant.scala 16:37]
  assign quant_unit_7_io_scale = io_scale; // @[quant.scala 17:32]
  assign quant_unit_7_io_shift = io_shift; // @[quant.scala 18:32]
  assign quant_unit_7_io_zero_point = io_zero_point; // @[quant.scala 19:37]
endmodule
module yolov8_maxpool_data_rwcontrol(
  input         clock,
  input         reset,
  input         io_pool_enable,
  input  [7:0]  io_zero_point,
  output        io_pool_finish,
  output [7:0]  io_pool_input_0,
  output [7:0]  io_pool_input_1,
  output [7:0]  io_pool_input_2,
  output [7:0]  io_pool_input_3,
  output [7:0]  io_pool_input_4,
  output [7:0]  io_pool_input_5,
  output [7:0]  io_pool_input_6,
  output [7:0]  io_pool_input_7,
  output        io_last_data_of_row,
  input         io_pool_outdata_valid,
  output [11:0] io_ofm_write_addr,
  output        io_ofm_en_write,
  output [11:0] io_ofm_read_addr,
  input  [63:0] io_ofm_read_bundle,
  input  [9:0]  io_row,
  input  [9:0]  io_col
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pool_cnt; // @[pool.scala 32:27]
  reg [1:0] pool_cnt_write; // @[pool.scala 34:31]
  reg  pool_enable_upedge_REG; // @[utils.scala 10:17]
  wire  pool_enable_upedge = ~pool_enable_upedge_REG & io_pool_enable; // @[utils.scala 10:27]
  reg [1:0] state; // @[pool.scala 39:22]
  reg [9:0] row_cnt; // @[pool.scala 106:30]
  wire [9:0] _pool_finish_once_T_1 = io_row - 10'h1; // @[pool.scala 114:45]
  wire [3:0] _pool_finish_once_T_2 = 2'h2 * 2'h2; // @[pool.scala 114:53]
  wire [9:0] _GEN_18 = {{6'd0}, _pool_finish_once_T_2}; // @[pool.scala 114:49]
  wire [9:0] _pool_finish_once_T_4 = _pool_finish_once_T_1 + _GEN_18; // @[pool.scala 114:49]
  reg [9:0] col_cnt; // @[pool.scala 107:30]
  wire [9:0] _last_data_of_row_T_1 = io_col - 10'h1; // @[pool.scala 113:49]
  wire [9:0] _last_data_of_row_T_4 = _last_data_of_row_T_1 + _GEN_18; // @[pool.scala 113:53]
  wire  last_data_of_row = col_cnt == _last_data_of_row_T_4; // @[pool.scala 113:38]
  wire  pool_finish_once = row_cnt == _pool_finish_once_T_4 & last_data_of_row; // @[pool.scala 114:62]
  wire [1:0] _pool_cnt_T_1 = pool_cnt + 2'h1; // @[pool.scala 60:37]
  wire [1:0] _GEN_2 = pool_cnt == 2'h2 ? 2'h0 : _pool_cnt_T_1; // @[pool.scala 56:47 57:26 60:26]
  wire [1:0] _GEN_3 = pool_cnt == 2'h2 ? 2'h2 : 2'h1; // @[pool.scala 56:47 58:22 61:22]
  reg [11:0] ofm_offset_write_addr; // @[pool.scala 101:40]
  wire  _write_last_data_T = ofm_offset_write_addr == 12'h18f; // @[pool.scala 149:44]
  reg [9:0] write_row_cnt; // @[pool.scala 129:36]
  wire  ofm_en_write = io_pool_outdata_valid & write_row_cnt >= 10'h4; // @[pool.scala 135:47]
  wire  write_last_data = ofm_offset_write_addr == 12'h18f & ofm_en_write; // @[pool.scala 149:89]
  wire [1:0] _GEN_4 = write_last_data ? 2'h0 : 2'h2; // @[pool.scala 65:34 66:22 68:22]
  wire [1:0] _GEN_5 = 2'h2 == state ? _GEN_4 : state; // @[pool.scala 40:18 39:22]
  wire  state_is_idle = state == 2'h0; // @[pool.scala 72:29]
  wire  state_is_pool = state == 2'h1; // @[pool.scala 73:29]
  wire  state_is_pool_finish_once = state == 2'h3; // @[pool.scala 74:41]
  wire  state_is_all_finish = state == 2'h2; // @[pool.scala 75:35]
  reg [11:0] ofm_base_read_addr; // @[pool.scala 78:37]
  reg [11:0] ofm_base_write_addr; // @[pool.scala 79:38]
  wire [10:0] _ofm_base_read_addr_T = pool_cnt * 9'h190; // @[pool.scala 80:33]
  wire [10:0] _ofm_base_write_addr_T = pool_cnt_write * 9'h190; // @[pool.scala 82:40]
  reg  zero_enable_reg; // @[pool.scala 108:38]
  wire [63:0] pool_in_data = zero_enable_reg ? {{56'd0}, io_zero_point} : io_ofm_read_bundle; // @[pool.scala 140:28]
  wire  clr_pool = reset | state_is_idle | state_is_pool_finish_once; // @[pool.scala 104:49]
  wire [9:0] _zero_enable_wire_T_4 = io_row + 10'h2; // @[pool.scala 110:89]
  wire [9:0] _zero_enable_wire_T_6 = _zero_enable_wire_T_4 - 10'h1; // @[pool.scala 110:97]
  wire [9:0] _zero_enable_wire_T_10 = io_col + 10'h2; // @[pool.scala 110:125]
  wire [9:0] _zero_enable_wire_T_12 = _zero_enable_wire_T_10 - 10'h1; // @[pool.scala 110:133]
  wire  zero_enable_wire = row_cnt < 10'h2 | col_cnt < 10'h2 | row_cnt > _zero_enable_wire_T_6 | col_cnt >
    _zero_enable_wire_T_12; // @[pool.scala 110:104]
  reg [11:0] ofm_offset_read_addr; // @[pool.scala 116:43]
  wire [9:0] _row_cnt_T_1 = row_cnt + 10'h1; // @[pool.scala 120:33]
  wire [9:0] _col_cnt_T_1 = col_cnt + 10'h1; // @[pool.scala 122:33]
  wire [11:0] _ofm_offset_read_addr_T_1 = ofm_offset_read_addr + 12'h1; // @[pool.scala 126:57]
  reg [9:0] write_col_cnt; // @[pool.scala 130:36]
  wire  _write_col_cnt_T = write_col_cnt == 10'h13; // @[pool.scala 131:67]
  wire [9:0] _write_col_cnt_T_2 = write_col_cnt + 10'h1; // @[pool.scala 131:92]
  wire [9:0] _write_row_cnt_T_2 = write_row_cnt + 10'h1; // @[pool.scala 132:88]
  reg  io_last_data_of_row_REG; // @[pool.scala 142:37]
  wire [1:0] _pool_cnt_write_T_1 = pool_cnt_write + 2'h1; // @[pool.scala 144:83]
  wire [11:0] _ofm_offset_write_addr_T_2 = ofm_offset_write_addr + 12'h1; // @[pool.scala 147:128]
  reg  io_pool_finish_REG; // @[utils.scala 19:16]
  assign io_pool_finish = io_pool_finish_REG & ~state_is_all_finish; // @[utils.scala 19:26]
  assign io_pool_input_0 = pool_in_data[7:0]; // @[pool.scala 94:38]
  assign io_pool_input_1 = pool_in_data[15:8]; // @[pool.scala 94:38]
  assign io_pool_input_2 = pool_in_data[23:16]; // @[pool.scala 94:38]
  assign io_pool_input_3 = pool_in_data[31:24]; // @[pool.scala 94:38]
  assign io_pool_input_4 = pool_in_data[39:32]; // @[pool.scala 94:38]
  assign io_pool_input_5 = pool_in_data[47:40]; // @[pool.scala 94:38]
  assign io_pool_input_6 = pool_in_data[55:48]; // @[pool.scala 94:38]
  assign io_pool_input_7 = pool_in_data[63:56]; // @[pool.scala 94:38]
  assign io_last_data_of_row = io_last_data_of_row_REG; // @[pool.scala 142:28]
  assign io_ofm_write_addr = ofm_base_write_addr + ofm_offset_write_addr; // @[pool.scala 138:47]
  assign io_ofm_en_write = io_pool_outdata_valid & write_row_cnt >= 10'h4; // @[pool.scala 135:47]
  assign io_ofm_read_addr = ofm_base_read_addr + ofm_offset_read_addr; // @[pool.scala 137:45]
  always @(posedge clock) begin
    if (reset) begin // @[pool.scala 32:27]
      pool_cnt <= 2'h0; // @[pool.scala 32:27]
    end else if (!(2'h0 == state)) begin // @[pool.scala 40:18]
      if (!(2'h1 == state)) begin // @[pool.scala 40:18]
        if (2'h3 == state) begin // @[pool.scala 40:18]
          pool_cnt <= _GEN_2;
        end
      end
    end
    if (reset) begin // @[pool.scala 34:31]
      pool_cnt_write <= 2'h1; // @[pool.scala 34:31]
    end else if (state_is_all_finish) begin // @[pool.scala 144:24]
      pool_cnt_write <= 2'h1;
    end else if (write_last_data) begin // @[pool.scala 144:52]
      pool_cnt_write <= _pool_cnt_write_T_1;
    end
    if (reset) begin // @[utils.scala 10:17]
      pool_enable_upedge_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      pool_enable_upedge_REG <= io_pool_enable; // @[utils.scala 10:17]
    end
    if (reset) begin // @[pool.scala 39:22]
      state <= 2'h0; // @[pool.scala 39:22]
    end else if (2'h0 == state) begin // @[pool.scala 40:18]
      if (pool_enable_upedge) begin // @[pool.scala 42:37]
        state <= 2'h1; // @[pool.scala 43:23]
      end else begin
        state <= 2'h0; // @[pool.scala 45:23]
      end
    end else if (2'h1 == state) begin // @[pool.scala 40:18]
      if (pool_finish_once) begin // @[pool.scala 49:35]
        state <= 2'h3; // @[pool.scala 50:22]
      end else begin
        state <= 2'h1; // @[pool.scala 52:22]
      end
    end else if (2'h3 == state) begin // @[pool.scala 40:18]
      state <= _GEN_3;
    end else begin
      state <= _GEN_5;
    end
    if (clr_pool) begin // @[pool.scala 106:30]
      row_cnt <= 10'h0; // @[pool.scala 106:30]
    end else if (state_is_pool) begin // @[pool.scala 117:28]
      if (last_data_of_row) begin // @[pool.scala 118:51]
        row_cnt <= _row_cnt_T_1; // @[pool.scala 120:24]
      end
    end
    if (clr_pool) begin // @[pool.scala 107:30]
      col_cnt <= 10'h0; // @[pool.scala 107:30]
    end else if (state_is_pool) begin // @[pool.scala 117:28]
      if (last_data_of_row) begin // @[pool.scala 118:51]
        col_cnt <= 10'h0; // @[pool.scala 119:25]
      end else begin
        col_cnt <= _col_cnt_T_1; // @[pool.scala 122:24]
      end
    end
    if (reset) begin // @[pool.scala 101:40]
      ofm_offset_write_addr <= 12'h0; // @[pool.scala 101:40]
    end else if (ofm_en_write) begin // @[pool.scala 146:23]
      if (_write_last_data_T) begin // @[pool.scala 147:36]
        ofm_offset_write_addr <= 12'h0;
      end else begin
        ofm_offset_write_addr <= _ofm_offset_write_addr_T_2;
      end
    end
    if (clr_pool) begin // @[pool.scala 129:36]
      write_row_cnt <= 10'h0; // @[pool.scala 129:36]
    end else if (io_pool_outdata_valid) begin // @[pool.scala 132:27]
      if (_write_col_cnt_T) begin // @[pool.scala 132:53]
        write_row_cnt <= _write_row_cnt_T_2;
      end
    end
    if (reset) begin // @[pool.scala 78:37]
      ofm_base_read_addr <= 12'h0; // @[pool.scala 78:37]
    end else begin
      ofm_base_read_addr <= {{1'd0}, _ofm_base_read_addr_T}; // @[pool.scala 80:23]
    end
    if (reset) begin // @[pool.scala 79:38]
      ofm_base_write_addr <= 12'h0; // @[pool.scala 79:38]
    end else begin
      ofm_base_write_addr <= {{1'd0}, _ofm_base_write_addr_T}; // @[pool.scala 82:24]
    end
    if (clr_pool) begin // @[pool.scala 108:38]
      zero_enable_reg <= 1'h0; // @[pool.scala 108:38]
    end else begin
      zero_enable_reg <= zero_enable_wire; // @[pool.scala 111:24]
    end
    if (clr_pool) begin // @[pool.scala 116:43]
      ofm_offset_read_addr <= 12'h0; // @[pool.scala 116:43]
    end else if (state_is_pool & ~zero_enable_wire) begin // @[pool.scala 125:50]
      ofm_offset_read_addr <= _ofm_offset_read_addr_T_1; // @[pool.scala 126:34]
    end
    if (clr_pool) begin // @[pool.scala 130:36]
      write_col_cnt <= 10'h0; // @[pool.scala 130:36]
    end else if (io_pool_outdata_valid) begin // @[pool.scala 131:27]
      if (write_col_cnt == 10'h13) begin // @[pool.scala 131:53]
        write_col_cnt <= 10'h0;
      end else begin
        write_col_cnt <= _write_col_cnt_T_2;
      end
    end
    io_last_data_of_row_REG <= col_cnt == _last_data_of_row_T_4; // @[pool.scala 113:38]
    if (reset) begin // @[utils.scala 19:16]
      io_pool_finish_REG <= 1'h0; // @[utils.scala 19:16]
    end else begin
      io_pool_finish_REG <= state_is_all_finish; // @[utils.scala 19:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pool_cnt = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  pool_cnt_write = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  pool_enable_upedge_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  row_cnt = _RAND_4[9:0];
  _RAND_5 = {1{`RANDOM}};
  col_cnt = _RAND_5[9:0];
  _RAND_6 = {1{`RANDOM}};
  ofm_offset_write_addr = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  write_row_cnt = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  ofm_base_read_addr = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  ofm_base_write_addr = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  zero_enable_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ofm_offset_read_addr = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  write_col_cnt = _RAND_12[9:0];
  _RAND_13 = {1{`RANDOM}};
  io_last_data_of_row_REG = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  io_pool_finish_REG = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module compare2(
  input        clock,
  input        reset,
  input  [7:0] io_a,
  input  [7:0] io_b,
  output [7:0] io_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] out; // @[pool.scala 272:26]
  wire  valid = io_a < io_b; // @[pool.scala 275:27]
  assign io_dout = out; // @[pool.scala 277:16]
  always @(posedge clock) begin
    if (reset) begin // @[pool.scala 272:26]
      out <= 8'h0; // @[pool.scala 272:26]
    end else if (valid) begin // @[pool.scala 276:19]
      out <= io_b;
    end else begin
      out <= io_a;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cmp5(
  input        clock,
  input        reset,
  input  [7:0] io_in_0,
  input  [7:0] io_in_1,
  input  [7:0] io_in_2,
  input  [7:0] io_in_3,
  input  [7:0] io_in_4,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  cmp_0_clock; // @[pool.scala 244:33]
  wire  cmp_0_reset; // @[pool.scala 244:33]
  wire [7:0] cmp_0_io_a; // @[pool.scala 244:33]
  wire [7:0] cmp_0_io_b; // @[pool.scala 244:33]
  wire [7:0] cmp_0_io_dout; // @[pool.scala 244:33]
  wire  cmp_1_clock; // @[pool.scala 244:33]
  wire  cmp_1_reset; // @[pool.scala 244:33]
  wire [7:0] cmp_1_io_a; // @[pool.scala 244:33]
  wire [7:0] cmp_1_io_b; // @[pool.scala 244:33]
  wire [7:0] cmp_1_io_dout; // @[pool.scala 244:33]
  wire  cmp_2_clock; // @[pool.scala 244:33]
  wire  cmp_2_reset; // @[pool.scala 244:33]
  wire [7:0] cmp_2_io_a; // @[pool.scala 244:33]
  wire [7:0] cmp_2_io_b; // @[pool.scala 244:33]
  wire [7:0] cmp_2_io_dout; // @[pool.scala 244:33]
  wire  cmp_3_clock; // @[pool.scala 244:33]
  wire  cmp_3_reset; // @[pool.scala 244:33]
  wire [7:0] cmp_3_io_a; // @[pool.scala 244:33]
  wire [7:0] cmp_3_io_b; // @[pool.scala 244:33]
  wire [7:0] cmp_3_io_dout; // @[pool.scala 244:33]
  reg [7:0] temp_0; // @[pool.scala 241:25]
  reg [7:0] temp; // @[pool.scala 242:23]
  compare2 cmp_0 ( // @[pool.scala 244:33]
    .clock(cmp_0_clock),
    .reset(cmp_0_reset),
    .io_a(cmp_0_io_a),
    .io_b(cmp_0_io_b),
    .io_dout(cmp_0_io_dout)
  );
  compare2 cmp_1 ( // @[pool.scala 244:33]
    .clock(cmp_1_clock),
    .reset(cmp_1_reset),
    .io_a(cmp_1_io_a),
    .io_b(cmp_1_io_b),
    .io_dout(cmp_1_io_dout)
  );
  compare2 cmp_2 ( // @[pool.scala 244:33]
    .clock(cmp_2_clock),
    .reset(cmp_2_reset),
    .io_a(cmp_2_io_a),
    .io_b(cmp_2_io_b),
    .io_dout(cmp_2_io_dout)
  );
  compare2 cmp_3 ( // @[pool.scala 244:33]
    .clock(cmp_3_clock),
    .reset(cmp_3_reset),
    .io_a(cmp_3_io_a),
    .io_b(cmp_3_io_b),
    .io_dout(cmp_3_io_dout)
  );
  assign io_out = cmp_3_io_dout; // @[pool.scala 253:12]
  assign cmp_0_clock = clock;
  assign cmp_0_reset = reset;
  assign cmp_0_io_a = io_in_0; // @[pool.scala 245:17]
  assign cmp_0_io_b = io_in_1; // @[pool.scala 246:17]
  assign cmp_1_clock = clock;
  assign cmp_1_reset = reset;
  assign cmp_1_io_a = io_in_2; // @[pool.scala 247:17]
  assign cmp_1_io_b = io_in_3; // @[pool.scala 248:17]
  assign cmp_2_clock = clock;
  assign cmp_2_reset = reset;
  assign cmp_2_io_a = cmp_0_io_dout; // @[pool.scala 249:17]
  assign cmp_2_io_b = cmp_1_io_dout; // @[pool.scala 250:17]
  assign cmp_3_clock = clock;
  assign cmp_3_reset = reset;
  assign cmp_3_io_a = cmp_2_io_dout; // @[pool.scala 251:17]
  assign cmp_3_io_b = temp; // @[pool.scala 252:17]
  always @(posedge clock) begin
    temp_0 <= io_in_4; // @[pool.scala 241:25]
    temp <= temp_0; // @[pool.scala 242:23]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  temp = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pool_line_column(
  input        clock,
  input        reset,
  input  [7:0] io_input,
  input        io_pool_col_en,
  output [7:0] io_output
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
`endif // RANDOMIZE_REG_INIT
  wire  cmp_clock; // @[pool.scala 227:21]
  wire  cmp_reset; // @[pool.scala 227:21]
  wire [7:0] cmp_io_in_0; // @[pool.scala 227:21]
  wire [7:0] cmp_io_in_1; // @[pool.scala 227:21]
  wire [7:0] cmp_io_in_2; // @[pool.scala 227:21]
  wire [7:0] cmp_io_in_3; // @[pool.scala 227:21]
  wire [7:0] cmp_io_in_4; // @[pool.scala 227:21]
  wire [7:0] cmp_io_out; // @[pool.scala 227:21]
  reg [7:0] line_shift_1_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_1; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_2; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_3; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_4; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_5; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_6; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_7; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_8; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_9; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_10; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_11; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_12; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_13; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_14; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_15; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_16; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_17; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4_r_18; // @[Reg.scala 35:20]
  reg [7:0] line_shift_4; // @[Reg.scala 35:20]
  cmp5 cmp ( // @[pool.scala 227:21]
    .clock(cmp_clock),
    .reset(cmp_reset),
    .io_in_0(cmp_io_in_0),
    .io_in_1(cmp_io_in_1),
    .io_in_2(cmp_io_in_2),
    .io_in_3(cmp_io_in_3),
    .io_in_4(cmp_io_in_4),
    .io_out(cmp_io_out)
  );
  assign io_output = cmp_io_out; // @[pool.scala 233:15]
  assign cmp_clock = clock;
  assign cmp_reset = reset;
  assign cmp_io_in_0 = io_input; // @[pool.scala 228:18]
  assign cmp_io_in_1 = line_shift_1; // @[pool.scala 229:18]
  assign cmp_io_in_2 = line_shift_2; // @[pool.scala 230:18]
  assign cmp_io_in_3 = line_shift_3; // @[pool.scala 231:18]
  assign cmp_io_in_4 = line_shift_4; // @[pool.scala 232:18]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r <= io_input; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_1 <= line_shift_1_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_2 <= line_shift_1_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_3 <= line_shift_1_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_4 <= line_shift_1_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_5 <= line_shift_1_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_6 <= line_shift_1_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_7 <= line_shift_1_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_8 <= line_shift_1_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_9 <= line_shift_1_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_10 <= line_shift_1_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_11 <= line_shift_1_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_12 <= line_shift_1_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_13 <= line_shift_1_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_14 <= line_shift_1_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_15 <= line_shift_1_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_16 <= line_shift_1_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_17 <= line_shift_1_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1_r_18 <= line_shift_1_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_1 <= line_shift_1_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r <= line_shift_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_1 <= line_shift_2_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_2 <= line_shift_2_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_3 <= line_shift_2_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_4 <= line_shift_2_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_5 <= line_shift_2_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_6 <= line_shift_2_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_7 <= line_shift_2_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_8 <= line_shift_2_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_9 <= line_shift_2_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_10 <= line_shift_2_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_11 <= line_shift_2_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_12 <= line_shift_2_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_13 <= line_shift_2_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_14 <= line_shift_2_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_15 <= line_shift_2_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_16 <= line_shift_2_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_17 <= line_shift_2_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2_r_18 <= line_shift_2_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_2 <= line_shift_2_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r <= line_shift_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_1 <= line_shift_3_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_2 <= line_shift_3_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_3 <= line_shift_3_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_4 <= line_shift_3_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_5 <= line_shift_3_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_6 <= line_shift_3_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_7 <= line_shift_3_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_8 <= line_shift_3_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_9 <= line_shift_3_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_10 <= line_shift_3_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_11 <= line_shift_3_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_12 <= line_shift_3_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_13 <= line_shift_3_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_14 <= line_shift_3_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_15 <= line_shift_3_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_16 <= line_shift_3_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_17 <= line_shift_3_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3_r_18 <= line_shift_3_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_3 <= line_shift_3_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r <= line_shift_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_1 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_1 <= line_shift_4_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_2 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_2 <= line_shift_4_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_3 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_3 <= line_shift_4_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_4 <= line_shift_4_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_5 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_5 <= line_shift_4_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_6 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_6 <= line_shift_4_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_7 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_7 <= line_shift_4_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_8 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_8 <= line_shift_4_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_9 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_9 <= line_shift_4_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_10 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_10 <= line_shift_4_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_11 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_11 <= line_shift_4_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_12 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_12 <= line_shift_4_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_13 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_13 <= line_shift_4_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_14 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_14 <= line_shift_4_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_15 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_15 <= line_shift_4_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_16 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_16 <= line_shift_4_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_17 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_17 <= line_shift_4_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4_r_18 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4_r_18 <= line_shift_4_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      line_shift_4 <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_pool_col_en) begin // @[Reg.scala 36:18]
      line_shift_4 <= line_shift_4_r_18; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  line_shift_1_r = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  line_shift_1_r_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  line_shift_1_r_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  line_shift_1_r_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  line_shift_1_r_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  line_shift_1_r_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  line_shift_1_r_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  line_shift_1_r_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  line_shift_1_r_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  line_shift_1_r_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  line_shift_1_r_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  line_shift_1_r_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  line_shift_1_r_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  line_shift_1_r_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  line_shift_1_r_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  line_shift_1_r_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  line_shift_1_r_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  line_shift_1_r_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  line_shift_1_r_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  line_shift_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  line_shift_2_r = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  line_shift_2_r_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  line_shift_2_r_2 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  line_shift_2_r_3 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  line_shift_2_r_4 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  line_shift_2_r_5 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  line_shift_2_r_6 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  line_shift_2_r_7 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  line_shift_2_r_8 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  line_shift_2_r_9 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  line_shift_2_r_10 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  line_shift_2_r_11 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  line_shift_2_r_12 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  line_shift_2_r_13 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  line_shift_2_r_14 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  line_shift_2_r_15 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  line_shift_2_r_16 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  line_shift_2_r_17 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  line_shift_2_r_18 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  line_shift_2 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  line_shift_3_r = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  line_shift_3_r_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  line_shift_3_r_2 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  line_shift_3_r_3 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  line_shift_3_r_4 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  line_shift_3_r_5 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  line_shift_3_r_6 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  line_shift_3_r_7 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  line_shift_3_r_8 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  line_shift_3_r_9 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  line_shift_3_r_10 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  line_shift_3_r_11 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  line_shift_3_r_12 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  line_shift_3_r_13 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  line_shift_3_r_14 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  line_shift_3_r_15 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  line_shift_3_r_16 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  line_shift_3_r_17 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  line_shift_3_r_18 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  line_shift_3 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  line_shift_4_r = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  line_shift_4_r_1 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  line_shift_4_r_2 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  line_shift_4_r_3 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  line_shift_4_r_4 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  line_shift_4_r_5 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  line_shift_4_r_6 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  line_shift_4_r_7 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  line_shift_4_r_8 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  line_shift_4_r_9 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  line_shift_4_r_10 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  line_shift_4_r_11 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  line_shift_4_r_12 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  line_shift_4_r_13 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  line_shift_4_r_14 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  line_shift_4_r_15 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  line_shift_4_r_16 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  line_shift_4_r_17 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  line_shift_4_r_18 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  line_shift_4 = _RAND_79[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module compare_line_unit(
  input        clock,
  input        reset,
  input  [7:0] io_input,
  input        io_last_data_of_row,
  output [7:0] io_output,
  output       io_outdata_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  cmp_clock; // @[pool.scala 202:21]
  wire  cmp_reset; // @[pool.scala 202:21]
  wire [7:0] cmp_io_in_0; // @[pool.scala 202:21]
  wire [7:0] cmp_io_in_1; // @[pool.scala 202:21]
  wire [7:0] cmp_io_in_2; // @[pool.scala 202:21]
  wire [7:0] cmp_io_in_3; // @[pool.scala 202:21]
  wire [7:0] cmp_io_in_4; // @[pool.scala 202:21]
  wire [7:0] cmp_io_out; // @[pool.scala 202:21]
  wire  pool_column_clock; // @[pool.scala 211:29]
  wire  pool_column_reset; // @[pool.scala 211:29]
  wire [7:0] pool_column_io_input; // @[pool.scala 211:29]
  wire  pool_column_io_pool_col_en; // @[pool.scala 211:29]
  wire [7:0] pool_column_io_output; // @[pool.scala 211:29]
  reg  start; // @[pool.scala 180:24]
  reg  last_up_REG; // @[utils.scala 10:17]
  wire  last_up = ~last_up_REG & io_last_data_of_row; // @[utils.scala 10:27]
  reg  last_r; // @[Reg.scala 35:20]
  reg  last; // @[Reg.scala 35:20]
  reg [2:0] cnt; // @[pool.scala 185:22]
  wire  _start_T_1 = cnt == 3'h4; // @[pool.scala 186:52]
  wire  _start_T_2 = cnt == 3'h4 ? 1'h0 : start; // @[pool.scala 186:47]
  wire [2:0] _cnt_T_2 = cnt + 3'h1; // @[pool.scala 187:49]
  reg  valid_delay1; // @[pool.scala 192:29]
  reg  valid_delay2; // @[pool.scala 193:29]
  reg  valid_delay3; // @[pool.scala 194:29]
  reg [7:0] temp_0; // @[pool.scala 197:35]
  reg [7:0] temp_1; // @[pool.scala 197:35]
  reg [7:0] temp_2; // @[pool.scala 197:35]
  reg [7:0] temp_3; // @[pool.scala 197:35]
  cmp5 cmp ( // @[pool.scala 202:21]
    .clock(cmp_clock),
    .reset(cmp_reset),
    .io_in_0(cmp_io_in_0),
    .io_in_1(cmp_io_in_1),
    .io_in_2(cmp_io_in_2),
    .io_in_3(cmp_io_in_3),
    .io_in_4(cmp_io_in_4),
    .io_out(cmp_io_out)
  );
  pool_line_column pool_column ( // @[pool.scala 211:29]
    .clock(pool_column_clock),
    .reset(pool_column_reset),
    .io_input(pool_column_io_input),
    .io_pool_col_en(pool_column_io_pool_col_en),
    .io_output(pool_column_io_output)
  );
  assign io_output = pool_column_io_output; // @[pool.scala 214:15]
  assign io_outdata_valid = valid_delay3; // @[pool.scala 195:21]
  assign cmp_clock = clock;
  assign cmp_reset = reset;
  assign cmp_io_in_0 = temp_0; // @[pool.scala 208:26]
  assign cmp_io_in_1 = temp_1; // @[pool.scala 208:26]
  assign cmp_io_in_2 = temp_2; // @[pool.scala 208:26]
  assign cmp_io_in_3 = temp_3; // @[pool.scala 208:26]
  assign cmp_io_in_4 = io_input; // @[pool.scala 205:26]
  assign pool_column_clock = clock;
  assign pool_column_reset = reset;
  assign pool_column_io_input = cmp_io_out; // @[pool.scala 212:26]
  assign pool_column_io_pool_col_en = cnt == 3'h0; // @[pool.scala 190:19]
  always @(posedge clock) begin
    if (reset) begin // @[pool.scala 180:24]
      start <= 1'h0; // @[pool.scala 180:24]
    end else begin
      start <= last | _start_T_2; // @[pool.scala 186:11]
    end
    if (reset) begin // @[utils.scala 10:17]
      last_up_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      last_up_REG <= io_last_data_of_row; // @[utils.scala 10:17]
    end
    if (reset) begin // @[Reg.scala 35:20]
      last_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      last_r <= last_up;
    end
    if (reset) begin // @[Reg.scala 35:20]
      last <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      last <= last_r;
    end
    if (reset) begin // @[pool.scala 185:22]
      cnt <= 3'h0; // @[pool.scala 185:22]
    end else if (start) begin // @[pool.scala 187:15]
      if (_start_T_1) begin // @[pool.scala 187:26]
        cnt <= 3'h0;
      end else begin
        cnt <= _cnt_T_2;
      end
    end
    valid_delay1 <= cnt == 3'h0; // @[pool.scala 190:19]
    valid_delay2 <= valid_delay1; // @[pool.scala 193:29]
    valid_delay3 <= valid_delay2; // @[pool.scala 194:29]
    if (reset) begin // @[pool.scala 197:35]
      temp_0 <= 8'h0; // @[pool.scala 197:35]
    end else begin
      temp_0 <= temp_1; // @[pool.scala 200:17]
    end
    if (reset) begin // @[pool.scala 197:35]
      temp_1 <= 8'h0; // @[pool.scala 197:35]
    end else begin
      temp_1 <= temp_2; // @[pool.scala 200:17]
    end
    if (reset) begin // @[pool.scala 197:35]
      temp_2 <= 8'h0; // @[pool.scala 197:35]
    end else begin
      temp_2 <= temp_3; // @[pool.scala 200:17]
    end
    if (reset) begin // @[pool.scala 197:35]
      temp_3 <= 8'h0; // @[pool.scala 197:35]
    end else begin
      temp_3 <= io_input; // @[pool.scala 198:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  start = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  last_up_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  last_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  last = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cnt = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  valid_delay1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_delay2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  valid_delay3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  temp_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  temp_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  temp_2 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  temp_3 = _RAND_11[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MaxPool(
  input        clock,
  input        reset,
  input  [7:0] io_input_0,
  input  [7:0] io_input_1,
  input  [7:0] io_input_2,
  input  [7:0] io_input_3,
  input  [7:0] io_input_4,
  input  [7:0] io_input_5,
  input  [7:0] io_input_6,
  input  [7:0] io_input_7,
  input        io_last_data_of_row,
  output [7:0] io_output_0,
  output [7:0] io_output_1,
  output [7:0] io_output_2,
  output [7:0] io_output_3,
  output [7:0] io_output_4,
  output [7:0] io_output_5,
  output [7:0] io_output_6,
  output [7:0] io_output_7,
  output       io_outdata_valid
);
  wire  pool_0_clock; // @[pool.scala 163:49]
  wire  pool_0_reset; // @[pool.scala 163:49]
  wire [7:0] pool_0_io_input; // @[pool.scala 163:49]
  wire  pool_0_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_0_io_output; // @[pool.scala 163:49]
  wire  pool_0_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_1_clock; // @[pool.scala 163:49]
  wire  pool_1_reset; // @[pool.scala 163:49]
  wire [7:0] pool_1_io_input; // @[pool.scala 163:49]
  wire  pool_1_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_1_io_output; // @[pool.scala 163:49]
  wire  pool_1_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_2_clock; // @[pool.scala 163:49]
  wire  pool_2_reset; // @[pool.scala 163:49]
  wire [7:0] pool_2_io_input; // @[pool.scala 163:49]
  wire  pool_2_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_2_io_output; // @[pool.scala 163:49]
  wire  pool_2_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_3_clock; // @[pool.scala 163:49]
  wire  pool_3_reset; // @[pool.scala 163:49]
  wire [7:0] pool_3_io_input; // @[pool.scala 163:49]
  wire  pool_3_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_3_io_output; // @[pool.scala 163:49]
  wire  pool_3_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_4_clock; // @[pool.scala 163:49]
  wire  pool_4_reset; // @[pool.scala 163:49]
  wire [7:0] pool_4_io_input; // @[pool.scala 163:49]
  wire  pool_4_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_4_io_output; // @[pool.scala 163:49]
  wire  pool_4_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_5_clock; // @[pool.scala 163:49]
  wire  pool_5_reset; // @[pool.scala 163:49]
  wire [7:0] pool_5_io_input; // @[pool.scala 163:49]
  wire  pool_5_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_5_io_output; // @[pool.scala 163:49]
  wire  pool_5_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_6_clock; // @[pool.scala 163:49]
  wire  pool_6_reset; // @[pool.scala 163:49]
  wire [7:0] pool_6_io_input; // @[pool.scala 163:49]
  wire  pool_6_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_6_io_output; // @[pool.scala 163:49]
  wire  pool_6_io_outdata_valid; // @[pool.scala 163:49]
  wire  pool_7_clock; // @[pool.scala 163:49]
  wire  pool_7_reset; // @[pool.scala 163:49]
  wire [7:0] pool_7_io_input; // @[pool.scala 163:49]
  wire  pool_7_io_last_data_of_row; // @[pool.scala 163:49]
  wire [7:0] pool_7_io_output; // @[pool.scala 163:49]
  wire  pool_7_io_outdata_valid; // @[pool.scala 163:49]
  compare_line_unit pool_0 ( // @[pool.scala 163:49]
    .clock(pool_0_clock),
    .reset(pool_0_reset),
    .io_input(pool_0_io_input),
    .io_last_data_of_row(pool_0_io_last_data_of_row),
    .io_output(pool_0_io_output),
    .io_outdata_valid(pool_0_io_outdata_valid)
  );
  compare_line_unit pool_1 ( // @[pool.scala 163:49]
    .clock(pool_1_clock),
    .reset(pool_1_reset),
    .io_input(pool_1_io_input),
    .io_last_data_of_row(pool_1_io_last_data_of_row),
    .io_output(pool_1_io_output),
    .io_outdata_valid(pool_1_io_outdata_valid)
  );
  compare_line_unit pool_2 ( // @[pool.scala 163:49]
    .clock(pool_2_clock),
    .reset(pool_2_reset),
    .io_input(pool_2_io_input),
    .io_last_data_of_row(pool_2_io_last_data_of_row),
    .io_output(pool_2_io_output),
    .io_outdata_valid(pool_2_io_outdata_valid)
  );
  compare_line_unit pool_3 ( // @[pool.scala 163:49]
    .clock(pool_3_clock),
    .reset(pool_3_reset),
    .io_input(pool_3_io_input),
    .io_last_data_of_row(pool_3_io_last_data_of_row),
    .io_output(pool_3_io_output),
    .io_outdata_valid(pool_3_io_outdata_valid)
  );
  compare_line_unit pool_4 ( // @[pool.scala 163:49]
    .clock(pool_4_clock),
    .reset(pool_4_reset),
    .io_input(pool_4_io_input),
    .io_last_data_of_row(pool_4_io_last_data_of_row),
    .io_output(pool_4_io_output),
    .io_outdata_valid(pool_4_io_outdata_valid)
  );
  compare_line_unit pool_5 ( // @[pool.scala 163:49]
    .clock(pool_5_clock),
    .reset(pool_5_reset),
    .io_input(pool_5_io_input),
    .io_last_data_of_row(pool_5_io_last_data_of_row),
    .io_output(pool_5_io_output),
    .io_outdata_valid(pool_5_io_outdata_valid)
  );
  compare_line_unit pool_6 ( // @[pool.scala 163:49]
    .clock(pool_6_clock),
    .reset(pool_6_reset),
    .io_input(pool_6_io_input),
    .io_last_data_of_row(pool_6_io_last_data_of_row),
    .io_output(pool_6_io_output),
    .io_outdata_valid(pool_6_io_outdata_valid)
  );
  compare_line_unit pool_7 ( // @[pool.scala 163:49]
    .clock(pool_7_clock),
    .reset(pool_7_reset),
    .io_input(pool_7_io_input),
    .io_last_data_of_row(pool_7_io_last_data_of_row),
    .io_output(pool_7_io_output),
    .io_outdata_valid(pool_7_io_outdata_valid)
  );
  assign io_output_0 = pool_0_io_output; // @[pool.scala 167:22]
  assign io_output_1 = pool_1_io_output; // @[pool.scala 167:22]
  assign io_output_2 = pool_2_io_output; // @[pool.scala 167:22]
  assign io_output_3 = pool_3_io_output; // @[pool.scala 167:22]
  assign io_output_4 = pool_4_io_output; // @[pool.scala 167:22]
  assign io_output_5 = pool_5_io_output; // @[pool.scala 167:22]
  assign io_output_6 = pool_6_io_output; // @[pool.scala 167:22]
  assign io_output_7 = pool_7_io_output; // @[pool.scala 167:22]
  assign io_outdata_valid = pool_0_io_outdata_valid; // @[pool.scala 169:21]
  assign pool_0_clock = clock;
  assign pool_0_reset = reset;
  assign pool_0_io_input = io_input_0; // @[pool.scala 165:26]
  assign pool_0_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_1_clock = clock;
  assign pool_1_reset = reset;
  assign pool_1_io_input = io_input_1; // @[pool.scala 165:26]
  assign pool_1_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_2_clock = clock;
  assign pool_2_reset = reset;
  assign pool_2_io_input = io_input_2; // @[pool.scala 165:26]
  assign pool_2_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_3_clock = clock;
  assign pool_3_reset = reset;
  assign pool_3_io_input = io_input_3; // @[pool.scala 165:26]
  assign pool_3_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_4_clock = clock;
  assign pool_4_reset = reset;
  assign pool_4_io_input = io_input_4; // @[pool.scala 165:26]
  assign pool_4_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_5_clock = clock;
  assign pool_5_reset = reset;
  assign pool_5_io_input = io_input_5; // @[pool.scala 165:26]
  assign pool_5_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_6_clock = clock;
  assign pool_6_reset = reset;
  assign pool_6_io_input = io_input_6; // @[pool.scala 165:26]
  assign pool_6_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
  assign pool_7_clock = clock;
  assign pool_7_reset = reset;
  assign pool_7_io_input = io_input_7; // @[pool.scala 165:26]
  assign pool_7_io_last_data_of_row = io_last_data_of_row; // @[pool.scala 166:37]
endmodule
module BottleNeck_add(
  input         clock,
  input         reset,
  output [10:0] io_ifm_read_addr,
  output        io_ifm_addr_read_sel,
  input  [7:0]  io_ifm_read_data_0,
  input  [7:0]  io_ifm_read_data_1,
  input  [7:0]  io_ifm_read_data_2,
  input  [7:0]  io_ifm_read_data_3,
  input  [7:0]  io_ifm_read_data_4,
  input  [7:0]  io_ifm_read_data_5,
  input  [7:0]  io_ifm_read_data_6,
  input  [7:0]  io_ifm_read_data_7,
  output [11:0] io_ofm_write_addr,
  output        io_ofm_en_write,
  output [11:0] io_ofm_read_addr,
  output [63:0] io_ofm_write_data,
  input  [63:0] io_ofm_read_data,
  input  [9:0]  io_col,
  input  [9:0]  io_row,
  input         io_bottleneck_add_enable,
  output        io_bottleneck_add_finish,
  output [7:0]  io_bn_add_in0_0,
  output [7:0]  io_bn_add_in0_1,
  output [7:0]  io_bn_add_in0_2,
  output [7:0]  io_bn_add_in0_3,
  output [7:0]  io_bn_add_in0_4,
  output [7:0]  io_bn_add_in0_5,
  output [7:0]  io_bn_add_in0_6,
  output [7:0]  io_bn_add_in0_7,
  output [7:0]  io_bn_add_in1_0,
  output [7:0]  io_bn_add_in1_1,
  output [7:0]  io_bn_add_in1_2,
  output [7:0]  io_bn_add_in1_3,
  output [7:0]  io_bn_add_in1_4,
  output [7:0]  io_bn_add_in1_5,
  output [7:0]  io_bn_add_in1_6,
  output [7:0]  io_bn_add_in1_7,
  input  [7:0]  io_bn_add_result_0,
  input  [7:0]  io_bn_add_result_1,
  input  [7:0]  io_bn_add_result_2,
  input  [7:0]  io_bn_add_result_3,
  input  [7:0]  io_bn_add_result_4,
  input  [7:0]  io_bn_add_result_5,
  input  [7:0]  io_bn_add_result_6,
  input  [7:0]  io_bn_add_result_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
`endif // RANDOMIZE_REG_INIT
  reg  bottleneck_add_enable_upegde_REG; // @[utils.scala 10:17]
  wire  bottleneck_add_enable_upegde = ~bottleneck_add_enable_upegde_REG & io_bottleneck_add_enable; // @[utils.scala 10:27]
  reg  bn_add_working; // @[ofmBuffer.scala 59:31]
  reg [9:0] col_cnt; // @[ofmBuffer.scala 61:24]
  reg [9:0] row_cnt; // @[ofmBuffer.scala 62:24]
  wire [9:0] _col_cnt_T_1 = io_col - 10'h1; // @[ofmBuffer.scala 63:54]
  wire  _col_cnt_T_2 = col_cnt == _col_cnt_T_1; // @[ofmBuffer.scala 63:44]
  wire [9:0] _col_cnt_T_4 = col_cnt + 10'h1; // @[ofmBuffer.scala 63:71]
  wire [9:0] _row_cnt_T_4 = row_cnt + 10'h1; // @[ofmBuffer.scala 64:67]
  wire [9:0] _bn_finish_T_1 = io_row - 10'h1; // @[ofmBuffer.scala 67:34]
  wire  bn_finish = row_cnt == _bn_finish_T_1 & _col_cnt_T_2; // @[ofmBuffer.scala 67:40]
  reg  current_is_singal_or_double; // @[ofmBuffer.scala 70:44]
  wire  _current_is_singal_or_double_T_3 = ~current_is_singal_or_double; // @[ofmBuffer.scala 71:80]
  wire  _current_is_singal_or_double_T_4 = _col_cnt_T_2 ? ~current_is_singal_or_double : current_is_singal_or_double; // @[ofmBuffer.scala 71:56]
  reg [10:0] ifm_read_addr_singal; // @[ofmBuffer.scala 76:37]
  reg [10:0] ifm_read_addr_double; // @[ofmBuffer.scala 77:37]
  wire [10:0] _ifm_read_addr_singal_T_1 = ifm_read_addr_singal + 11'h1; // @[ofmBuffer.scala 78:84]
  wire [10:0] _ifm_read_addr_double_T_1 = ifm_read_addr_double + 11'h1; // @[ofmBuffer.scala 79:89]
  wire [11:0] _ifm_read_addr_T = {1'h0,ifm_read_addr_singal}; // @[Cat.scala 33:92]
  wire [11:0] _ifm_read_addr_T_1 = {1'h1,ifm_read_addr_double}; // @[Cat.scala 33:92]
  wire [11:0] ifm_read_addr = _current_is_singal_or_double_T_3 ? _ifm_read_addr_T : _ifm_read_addr_T_1; // @[ofmBuffer.scala 80:28]
  reg [11:0] ofm_read_addr; // @[ofmBuffer.scala 85:32]
  reg [11:0] ofm_write_addr_r; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_2; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_3; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_4; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_5; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_6; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_7; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_8; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_9; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_10; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_11; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_12; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_13; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_14; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_r_15; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr; // @[Reg.scala 35:20]
  reg  ofm_en_write_r; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_1; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_2; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_3; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_4; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_5; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_6; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_7; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_8; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_9; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_10; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_11; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_12; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_13; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_14; // @[Reg.scala 35:20]
  reg  ofm_en_write_r_15; // @[Reg.scala 35:20]
  reg  ofm_en_write; // @[Reg.scala 35:20]
  wire [11:0] _ofm_read_addr_T_1 = ofm_read_addr + 12'h1; // @[ofmBuffer.scala 88:52]
  wire [55:0] _io_ofm_write_data_T_5 = {io_bn_add_result_6,io_bn_add_result_5,io_bn_add_result_4,io_bn_add_result_3,
    io_bn_add_result_2,io_bn_add_result_1,io_bn_add_result_0}; // @[Cat.scala 33:92]
  reg  bn_finish_upedge_REG; // @[utils.scala 10:17]
  wire  bn_finish_upedge = ~bn_finish_upedge_REG & bn_finish; // @[utils.scala 10:27]
  reg  bottleneck_finish_r; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_1; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_2; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_3; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_4; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_5; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_6; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_7; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_8; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_9; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_10; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_11; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_12; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_13; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_14; // @[Reg.scala 35:20]
  reg  bottleneck_finish_r_15; // @[Reg.scala 35:20]
  reg  bottleneck_finish; // @[Reg.scala 35:20]
  assign io_ifm_read_addr = ifm_read_addr[11:1]; // @[ofmBuffer.scala 81:38]
  assign io_ifm_addr_read_sel = ifm_read_addr[0]; // @[ofmBuffer.scala 82:42]
  assign io_ofm_write_addr = ofm_write_addr; // @[ofmBuffer.scala 90:22]
  assign io_ofm_en_write = ofm_en_write; // @[ofmBuffer.scala 89:20]
  assign io_ofm_read_addr = ofm_read_addr; // @[ofmBuffer.scala 91:21]
  assign io_ofm_write_data = {io_bn_add_result_7,_io_ofm_write_data_T_5}; // @[Cat.scala 33:92]
  assign io_bottleneck_add_finish = bottleneck_finish; // @[ofmBuffer.scala 112:29]
  assign io_bn_add_in0_0 = io_ifm_read_data_0; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_1 = io_ifm_read_data_1; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_2 = io_ifm_read_data_2; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_3 = io_ifm_read_data_3; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_4 = io_ifm_read_data_4; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_5 = io_ifm_read_data_5; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_6 = io_ifm_read_data_6; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in0_7 = io_ifm_read_data_7; // @[ofmBuffer.scala 93:33 94:23]
  assign io_bn_add_in1_0 = io_ofm_read_data[7:0]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_1 = io_ofm_read_data[15:8]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_2 = io_ofm_read_data[23:16]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_3 = io_ofm_read_data[31:24]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_4 = io_ofm_read_data[39:32]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_5 = io_ofm_read_data[47:40]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_6 = io_ofm_read_data[55:48]; // @[ofmBuffer.scala 100:47]
  assign io_bn_add_in1_7 = io_ofm_read_data[63:56]; // @[ofmBuffer.scala 100:47]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 10:17]
      bottleneck_add_enable_upegde_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      bottleneck_add_enable_upegde_REG <= io_bottleneck_add_enable; // @[utils.scala 10:17]
    end
    if (reset) begin // @[ofmBuffer.scala 59:31]
      bn_add_working <= 1'h0; // @[ofmBuffer.scala 59:31]
    end else if (bn_finish) begin // @[ofmBuffer.scala 68:24]
      bn_add_working <= 1'h0;
    end else begin
      bn_add_working <= bottleneck_add_enable_upegde | bn_add_working;
    end
    if (reset) begin // @[ofmBuffer.scala 61:24]
      col_cnt <= 10'h0; // @[ofmBuffer.scala 61:24]
    end else if (bn_add_working) begin // @[ofmBuffer.scala 63:17]
      if (col_cnt == _col_cnt_T_1) begin // @[ofmBuffer.scala 63:36]
        col_cnt <= 10'h0;
      end else begin
        col_cnt <= _col_cnt_T_4;
      end
    end else begin
      col_cnt <= 10'h0;
    end
    if (reset) begin // @[ofmBuffer.scala 62:24]
      row_cnt <= 10'h0; // @[ofmBuffer.scala 62:24]
    end else if (bn_add_working) begin // @[ofmBuffer.scala 64:17]
      if (_col_cnt_T_2) begin // @[ofmBuffer.scala 64:36]
        row_cnt <= _row_cnt_T_4;
      end
    end else begin
      row_cnt <= 10'h0;
    end
    if (reset) begin // @[ofmBuffer.scala 70:44]
      current_is_singal_or_double <= 1'h0; // @[ofmBuffer.scala 70:44]
    end else begin
      current_is_singal_or_double <= bn_add_working & _current_is_singal_or_double_T_4; // @[ofmBuffer.scala 71:32]
    end
    if (reset) begin // @[ofmBuffer.scala 76:37]
      ifm_read_addr_singal <= 11'h0; // @[ofmBuffer.scala 76:37]
    end else if (bn_add_working) begin // @[ofmBuffer.scala 78:30]
      if (_current_is_singal_or_double_T_3) begin // @[ofmBuffer.scala 78:49]
        ifm_read_addr_singal <= _ifm_read_addr_singal_T_1;
      end
    end else begin
      ifm_read_addr_singal <= 11'h0;
    end
    if (reset) begin // @[ofmBuffer.scala 77:37]
      ifm_read_addr_double <= 11'h0; // @[ofmBuffer.scala 77:37]
    end else if (bn_add_working) begin // @[ofmBuffer.scala 79:32]
      if (current_is_singal_or_double) begin // @[ofmBuffer.scala 79:52]
        ifm_read_addr_double <= _ifm_read_addr_double_T_1;
      end
    end else begin
      ifm_read_addr_double <= 11'h0;
    end
    if (reset) begin // @[ofmBuffer.scala 85:32]
      ofm_read_addr <= 12'h0; // @[ofmBuffer.scala 85:32]
    end else if (bn_add_working) begin // @[ofmBuffer.scala 88:23]
      ofm_read_addr <= _ofm_read_addr_T_1;
    end else begin
      ofm_read_addr <= 12'h0;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r <= ofm_read_addr;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_1 <= ofm_write_addr_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_2 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_2 <= ofm_write_addr_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_3 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_3 <= ofm_write_addr_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_4 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_4 <= ofm_write_addr_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_5 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_5 <= ofm_write_addr_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_6 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_6 <= ofm_write_addr_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_7 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_7 <= ofm_write_addr_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_8 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_8 <= ofm_write_addr_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_9 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_9 <= ofm_write_addr_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_10 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_10 <= ofm_write_addr_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_11 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_11 <= ofm_write_addr_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_12 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_12 <= ofm_write_addr_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_13 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_13 <= ofm_write_addr_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_14 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_14 <= ofm_write_addr_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_r_15 <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr_r_15 <= ofm_write_addr_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr <= 12'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_write_addr <= ofm_write_addr_r_15;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r <= bn_add_working;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_1 <= ofm_en_write_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_2 <= ofm_en_write_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_3 <= ofm_en_write_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_4 <= ofm_en_write_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_5 <= ofm_en_write_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_6 <= ofm_en_write_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_7 <= ofm_en_write_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_8 <= ofm_en_write_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_9 <= ofm_en_write_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_10 <= ofm_en_write_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_11 <= ofm_en_write_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_12 <= ofm_en_write_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_13 <= ofm_en_write_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_14 <= ofm_en_write_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write_r_15 <= ofm_en_write_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_en_write <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      ofm_en_write <= ofm_en_write_r_15;
    end
    if (reset) begin // @[utils.scala 10:17]
      bn_finish_upedge_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      bn_finish_upedge_REG <= bn_finish; // @[utils.scala 10:17]
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r <= bn_finish_upedge;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_1 <= bottleneck_finish_r;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_2 <= bottleneck_finish_r_1;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_3 <= bottleneck_finish_r_2;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_4 <= bottleneck_finish_r_3;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_5 <= bottleneck_finish_r_4;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_6 <= bottleneck_finish_r_5;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_7 <= bottleneck_finish_r_6;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_8 <= bottleneck_finish_r_7;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_9 <= bottleneck_finish_r_8;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_10 <= bottleneck_finish_r_9;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_11 <= bottleneck_finish_r_10;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_12 <= bottleneck_finish_r_11;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_13 <= bottleneck_finish_r_12;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_14 <= bottleneck_finish_r_13;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish_r_15 <= bottleneck_finish_r_14;
    end
    if (reset) begin // @[Reg.scala 35:20]
      bottleneck_finish <= 1'h0; // @[Reg.scala 35:20]
    end else begin
      bottleneck_finish <= bottleneck_finish_r_15;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bottleneck_add_enable_upegde_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bn_add_working = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  col_cnt = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  row_cnt = _RAND_3[9:0];
  _RAND_4 = {1{`RANDOM}};
  current_is_singal_or_double = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  ifm_read_addr_singal = _RAND_5[10:0];
  _RAND_6 = {1{`RANDOM}};
  ifm_read_addr_double = _RAND_6[10:0];
  _RAND_7 = {1{`RANDOM}};
  ofm_read_addr = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  ofm_write_addr_r = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  ofm_write_addr_r_1 = _RAND_9[11:0];
  _RAND_10 = {1{`RANDOM}};
  ofm_write_addr_r_2 = _RAND_10[11:0];
  _RAND_11 = {1{`RANDOM}};
  ofm_write_addr_r_3 = _RAND_11[11:0];
  _RAND_12 = {1{`RANDOM}};
  ofm_write_addr_r_4 = _RAND_12[11:0];
  _RAND_13 = {1{`RANDOM}};
  ofm_write_addr_r_5 = _RAND_13[11:0];
  _RAND_14 = {1{`RANDOM}};
  ofm_write_addr_r_6 = _RAND_14[11:0];
  _RAND_15 = {1{`RANDOM}};
  ofm_write_addr_r_7 = _RAND_15[11:0];
  _RAND_16 = {1{`RANDOM}};
  ofm_write_addr_r_8 = _RAND_16[11:0];
  _RAND_17 = {1{`RANDOM}};
  ofm_write_addr_r_9 = _RAND_17[11:0];
  _RAND_18 = {1{`RANDOM}};
  ofm_write_addr_r_10 = _RAND_18[11:0];
  _RAND_19 = {1{`RANDOM}};
  ofm_write_addr_r_11 = _RAND_19[11:0];
  _RAND_20 = {1{`RANDOM}};
  ofm_write_addr_r_12 = _RAND_20[11:0];
  _RAND_21 = {1{`RANDOM}};
  ofm_write_addr_r_13 = _RAND_21[11:0];
  _RAND_22 = {1{`RANDOM}};
  ofm_write_addr_r_14 = _RAND_22[11:0];
  _RAND_23 = {1{`RANDOM}};
  ofm_write_addr_r_15 = _RAND_23[11:0];
  _RAND_24 = {1{`RANDOM}};
  ofm_write_addr = _RAND_24[11:0];
  _RAND_25 = {1{`RANDOM}};
  ofm_en_write_r = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ofm_en_write_r_1 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ofm_en_write_r_2 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  ofm_en_write_r_3 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  ofm_en_write_r_4 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  ofm_en_write_r_5 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  ofm_en_write_r_6 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  ofm_en_write_r_7 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  ofm_en_write_r_8 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  ofm_en_write_r_9 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ofm_en_write_r_10 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  ofm_en_write_r_11 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ofm_en_write_r_12 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ofm_en_write_r_13 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  ofm_en_write_r_14 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  ofm_en_write_r_15 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ofm_en_write = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  bn_finish_upedge_REG = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  bottleneck_finish_r = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  bottleneck_finish_r_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  bottleneck_finish_r_2 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  bottleneck_finish_r_3 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  bottleneck_finish_r_4 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  bottleneck_finish_r_5 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  bottleneck_finish_r_6 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  bottleneck_finish_r_7 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  bottleneck_finish_r_8 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  bottleneck_finish_r_9 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  bottleneck_finish_r_10 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  bottleneck_finish_r_11 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  bottleneck_finish_r_12 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  bottleneck_finish_r_13 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  bottleneck_finish_r_14 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  bottleneck_finish_r_15 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  bottleneck_finish = _RAND_59[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TPRAM_WRAP_96(
  input         clock,
  input         io_wen,
  input  [11:0] io_waddr,
  input  [11:0] io_raddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata
);
  wire  tpram_CLKA; // @[utils.scala 218:23]
  wire  tpram_CLKB; // @[utils.scala 218:23]
  wire  tpram_CENB; // @[utils.scala 218:23]
  wire  tpram_CENA; // @[utils.scala 218:23]
  wire [11:0] tpram_AB; // @[utils.scala 218:23]
  wire [11:0] tpram_AA; // @[utils.scala 218:23]
  wire [63:0] tpram_DB; // @[utils.scala 218:23]
  wire [63:0] tpram_QA; // @[utils.scala 218:23]
  TPRAM #(.DATA_WIDTH(64), .DEPTH(4096), .RAM_STYLE_VAL("block")) tpram ( // @[utils.scala 218:23]
    .CLKA(tpram_CLKA),
    .CLKB(tpram_CLKB),
    .CENB(tpram_CENB),
    .CENA(tpram_CENA),
    .AB(tpram_AB),
    .AA(tpram_AA),
    .DB(tpram_DB),
    .QA(tpram_QA)
  );
  assign io_rdata = tpram_QA; // @[utils.scala 230:12]
  assign tpram_CLKA = clock; // @[utils.scala 222:19]
  assign tpram_CLKB = clock; // @[utils.scala 223:19]
  assign tpram_CENB = ~io_wen; // @[utils.scala 224:22]
  assign tpram_CENA = 1'h0; // @[utils.scala 225:22]
  assign tpram_AB = io_waddr; // @[utils.scala 226:17]
  assign tpram_AA = io_raddr; // @[utils.scala 227:17]
  assign tpram_DB = io_wdata; // @[utils.scala 228:17]
endmodule
module OfmBuffer(
  input         clock,
  input  [11:0] io_bram_write_addr,
  input         io_bram_en_write,
  input  [11:0] io_bram_read_addr,
  input  [63:0] io_ofm_store_bundle,
  output [63:0] io_ofm_out_bundle
);
  wire  TPRAM_WRAP_clock; // @[utils.scala 237:100]
  wire  TPRAM_WRAP_io_wen; // @[utils.scala 237:100]
  wire [11:0] TPRAM_WRAP_io_waddr; // @[utils.scala 237:100]
  wire [11:0] TPRAM_WRAP_io_raddr; // @[utils.scala 237:100]
  wire [63:0] TPRAM_WRAP_io_wdata; // @[utils.scala 237:100]
  wire [63:0] TPRAM_WRAP_io_rdata; // @[utils.scala 237:100]
  TPRAM_WRAP_96 TPRAM_WRAP ( // @[utils.scala 237:100]
    .clock(TPRAM_WRAP_clock),
    .io_wen(TPRAM_WRAP_io_wen),
    .io_waddr(TPRAM_WRAP_io_waddr),
    .io_raddr(TPRAM_WRAP_io_raddr),
    .io_wdata(TPRAM_WRAP_io_wdata),
    .io_rdata(TPRAM_WRAP_io_rdata)
  );
  assign io_ofm_out_bundle = TPRAM_WRAP_io_rdata; // @[ofmBuffer.scala 22:23]
  assign TPRAM_WRAP_clock = clock;
  assign TPRAM_WRAP_io_wen = io_bram_en_write; // @[ofmBuffer.scala 17:13]
  assign TPRAM_WRAP_io_waddr = io_bram_write_addr; // @[ofmBuffer.scala 19:15]
  assign TPRAM_WRAP_io_raddr = io_bram_read_addr; // @[ofmBuffer.scala 20:15]
  assign TPRAM_WRAP_io_wdata = io_ofm_store_bundle; // @[ofmBuffer.scala 21:15]
endmodule
module accel_top(
  input         clock,
  input         reset,
  input  [2:0]  io_sel,
  input  [10:0] io_ifmbuf_bram_addr_read_s1,
  input         io_ifmbuf_bram_addr_read_sel_s1,
  input  [9:0]  io_ifmbuf_bram_addr_read_s2_singal,
  input  [9:0]  io_ifmbuf_bram_addr_read_s2_double,
  input         io_ifmbuf_sel,
  input         io_ifmbuf_bram_en_write,
  input         io_recv_done,
  input         io_weightbuf_waddr_clear,
  input         io_weightbuf_bram_en_write,
  input  [6:0]  io_weightbuf_read_addr,
  input         io_kernal,
  input  [2:0]  io_weight_sel,
  input         io_biasbuf_waddr_clear,
  input         io_biasbuf_bram_en_write,
  input  [6:0]  io_biasbuf_read_addr,
  input         io_acc_read_en,
  input         io_acc_write_en,
  input  [11:0] io_acc_read_addr,
  input  [11:0] io_acc_write_addr,
  input         io_acc_prev_data_zero,
  input         io_acc_curr_data_zero,
  input         io_ofmbuf_bram_en_write,
  input  [11:0] io_ofmbuf_bram_write_addr,
  input  [63:0] io_ofmbuf_bram_read_addr,
  input  [9:0]  io_col,
  input  [9:0]  io_row,
  input         io_pad_top,
  input         io_pad_bottom,
  input         io_pad_left_and_right,
  input  [4:0]  io_zero_pad_valid_s2,
  input         io_zero_pad_valid_s1,
  input  [15:0] io_scale,
  input  [3:0]  io_shift,
  input  [7:0]  io_zero_point_in,
  input  [7:0]  io_zero_point_out,
  input  [7:0]  io_zero_point_A_act,
  input  [7:0]  io_ifm_in_0,
  input  [7:0]  io_ifm_in_1,
  input  [7:0]  io_ifm_in_2,
  input  [7:0]  io_ifm_in_3,
  input  [7:0]  io_ifm_in_4,
  input  [7:0]  io_ifm_in_5,
  input  [7:0]  io_ifm_in_6,
  input  [7:0]  io_ifm_in_7,
  input  [7:0]  io_weight_in_0,
  input  [7:0]  io_weight_in_1,
  input  [7:0]  io_weight_in_2,
  input  [7:0]  io_weight_in_3,
  input  [7:0]  io_weight_in_4,
  input  [7:0]  io_weight_in_5,
  input  [7:0]  io_weight_in_6,
  input  [7:0]  io_weight_in_7,
  input  [17:0] io_bias_in,
  input         io_bias_valid,
  output [63:0] io_ofm_out_bundle,
  input         io_skip_act,
  input         io_pool_enable,
  output        io_pool_finish,
  input         io_upsample_enable,
  input         io_bottleneck_add_enable,
  output        io_bottleneck_add_finish,
  input         io_s_mod,
  output [7:0]  io_act_indata_0,
  output [7:0]  io_act_indata_1,
  output [7:0]  io_act_indata_2,
  output [7:0]  io_act_indata_3,
  output [7:0]  io_act_indata_4,
  output [7:0]  io_act_indata_5,
  output [7:0]  io_act_indata_6,
  output [7:0]  io_act_indata_7,
  input  [7:0]  io_act_outdata_0,
  input  [7:0]  io_act_outdata_1,
  input  [7:0]  io_act_outdata_2,
  input  [7:0]  io_act_outdata_3,
  input  [7:0]  io_act_outdata_4,
  input  [7:0]  io_act_outdata_5,
  input  [7:0]  io_act_outdata_6,
  input  [7:0]  io_act_outdata_7,
  output [7:0]  io_bn_add_in0_0,
  output [7:0]  io_bn_add_in0_1,
  output [7:0]  io_bn_add_in0_2,
  output [7:0]  io_bn_add_in0_3,
  output [7:0]  io_bn_add_in0_4,
  output [7:0]  io_bn_add_in0_5,
  output [7:0]  io_bn_add_in0_6,
  output [7:0]  io_bn_add_in0_7,
  output [7:0]  io_bn_add_in1_0,
  output [7:0]  io_bn_add_in1_1,
  output [7:0]  io_bn_add_in1_2,
  output [7:0]  io_bn_add_in1_3,
  output [7:0]  io_bn_add_in1_4,
  output [7:0]  io_bn_add_in1_5,
  output [7:0]  io_bn_add_in1_6,
  output [7:0]  io_bn_add_in1_7,
  input  [7:0]  io_bn_add_result_0,
  input  [7:0]  io_bn_add_result_1,
  input  [7:0]  io_bn_add_result_2,
  input  [7:0]  io_bn_add_result_3,
  input  [7:0]  io_bn_add_result_4,
  input  [7:0]  io_bn_add_result_5,
  input  [7:0]  io_bn_add_result_6,
  input  [7:0]  io_bn_add_result_7,
  input         io_yolo_cls_en,
  output [63:0] io_yolo_cls_data_before_compare,
  input  [63:0] io_yolo_cls_data_after_compare
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  ifm_buf_clock; // @[acccel_top.scala 95:25]
  wire  ifm_buf_reset; // @[acccel_top.scala 95:25]
  wire [10:0] ifm_buf_io_ifmbuf_bram_addr_read_s1; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_ifmbuf_bram_addr_read_sel_s1; // @[acccel_top.scala 95:25]
  wire [9:0] ifm_buf_io_ifmbuf_bram_addr_read_s2_singal; // @[acccel_top.scala 95:25]
  wire [9:0] ifm_buf_io_ifmbuf_bram_addr_read_s2_double; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_bram_en_write; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_upsample_enable; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_recv_done; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_buf_sel; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_s_mod; // @[acccel_top.scala 95:25]
  wire [9:0] ifm_buf_io_col; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_0; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_1; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_2; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_3; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_4; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_5; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_6; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_in_7; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_0; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_1; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_2; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_3; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_4; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_5; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_6; // @[acccel_top.scala 95:25]
  wire [31:0] ifm_buf_io_ifm_o_data_7; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_pad_top; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_pad_bottom; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_pad_left_and_right; // @[acccel_top.scala 95:25]
  wire [4:0] ifm_buf_io_zero_pad_valid_s2; // @[acccel_top.scala 95:25]
  wire  ifm_buf_io_zero_pad_valid_s1; // @[acccel_top.scala 95:25]
  wire [7:0] ifm_buf_io_zero_point_in; // @[acccel_top.scala 95:25]
  wire  weight_buf_clock; // @[acccel_top.scala 120:28]
  wire  weight_buf_reset; // @[acccel_top.scala 120:28]
  wire  weight_buf_io_clear; // @[acccel_top.scala 120:28]
  wire  weight_buf_io_bram_write_en; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_0; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_1; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_2; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_3; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_4; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_5; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_6; // @[acccel_top.scala 120:28]
  wire [7:0] weight_buf_io_in_7; // @[acccel_top.scala 120:28]
  wire [6:0] weight_buf_io_read_addr; // @[acccel_top.scala 120:28]
  wire [2:0] weight_buf_io_sel_when_kernal_is_1; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_0; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_1; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_2; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_3; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_4; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_5; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_6; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_7; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_8; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_9; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_10; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_11; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_12; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_13; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_14; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_15; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_16; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_17; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_18; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_19; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_20; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_21; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_22; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_23; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_24; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_25; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_26; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_27; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_28; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_29; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_30; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_31; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_32; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_33; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_34; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_35; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_36; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_37; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_38; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_39; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_40; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_41; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_42; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_43; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_44; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_45; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_46; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_47; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_48; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_49; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_50; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_51; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_52; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_53; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_54; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_55; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_56; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_57; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_58; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_59; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_60; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_61; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_62; // @[acccel_top.scala 120:28]
  wire [71:0] weight_buf_io_weight_out_63; // @[acccel_top.scala 120:28]
  wire  weight_buf_io_kernal; // @[acccel_top.scala 120:28]
  wire  bias_buf_clock; // @[acccel_top.scala 134:26]
  wire  bias_buf_reset; // @[acccel_top.scala 134:26]
  wire  bias_buf_io_clear; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_in; // @[acccel_top.scala 134:26]
  wire [6:0] bias_buf_io_bram_addr_read; // @[acccel_top.scala 134:26]
  wire  bias_buf_io_bram_en_write; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_0; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_1; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_2; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_3; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_4; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_5; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_6; // @[acccel_top.scala 134:26]
  wire [17:0] bias_buf_io_bias_data_7; // @[acccel_top.scala 134:26]
  wire  sub_zero_clock; // @[acccel_top.scala 144:26]
  wire  sub_zero_reset; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_zero_point; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_0; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_1; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_2; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_3; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_4; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_5; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_6; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_7; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_8; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_9; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_10; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_11; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_12; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_13; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_14; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_15; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_16; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_17; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_18; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_19; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_20; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_21; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_22; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_23; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_24; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_25; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_26; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_27; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_28; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_29; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_30; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_in_31; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_0; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_1; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_2; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_3; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_4; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_5; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_6; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_7; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_8; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_9; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_10; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_11; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_12; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_13; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_14; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_15; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_16; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_17; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_18; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_19; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_20; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_21; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_22; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_23; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_24; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_25; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_26; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_27; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_28; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_29; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_30; // @[acccel_top.scala 144:26]
  wire [7:0] sub_zero_io_data_out_31; // @[acccel_top.scala 144:26]
  wire  line_buf_clock; // @[acccel_top.scala 154:26]
  wire  line_buf_reset; // @[acccel_top.scala 154:26]
  wire [2:0] line_buf_io_sel; // @[acccel_top.scala 154:26]
  wire  line_buf_io_s_mod; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_0; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_1; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_2; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_3; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_4; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_5; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_6; // @[acccel_top.scala 154:26]
  wire [31:0] line_buf_io_lineBuffer_i_data_7; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_0; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_1; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_2; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_3; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_4; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_5; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_6; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_7; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_8; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_9; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_10; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_11; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_12; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_13; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_14; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_15; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_16; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_17; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_18; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_19; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_20; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_21; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_22; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_23; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_24; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_25; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_26; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_27; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_28; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_29; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_30; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_31; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_32; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_33; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_34; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_35; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_36; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_37; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_38; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_39; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_40; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_41; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_42; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_43; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_44; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_45; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_46; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_47; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_48; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_49; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_50; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_51; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_52; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_53; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_54; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_55; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_56; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_57; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_58; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_59; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_60; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_61; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_62; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_63; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_64; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_65; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_66; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_67; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_68; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_69; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_70; // @[acccel_top.scala 154:26]
  wire [7:0] line_buf_io_lineBuffer_o_data_71; // @[acccel_top.scala 154:26]
  wire  conv_clock; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_0; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_1; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_2; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_3; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_4; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_5; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_6; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_7; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_8; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_9; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_10; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_11; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_12; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_13; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_14; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_15; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_16; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_17; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_18; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_19; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_20; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_21; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_22; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_23; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_24; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_25; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_26; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_27; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_28; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_29; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_30; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_31; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_32; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_33; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_34; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_35; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_36; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_37; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_38; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_39; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_40; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_41; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_42; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_43; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_44; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_45; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_46; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_47; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_48; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_49; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_50; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_51; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_52; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_53; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_54; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_55; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_56; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_57; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_58; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_59; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_60; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_61; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_62; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_63; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_64; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_65; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_66; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_67; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_68; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_69; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_70; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_ifm_win_33_71; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_0; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_1; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_2; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_3; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_4; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_5; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_6; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_7; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_8; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_9; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_10; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_11; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_12; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_13; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_14; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_15; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_16; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_17; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_18; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_19; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_20; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_21; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_22; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_23; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_24; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_25; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_26; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_27; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_28; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_29; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_30; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_31; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_32; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_33; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_34; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_35; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_36; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_37; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_38; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_39; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_40; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_41; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_42; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_43; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_44; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_45; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_46; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_47; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_48; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_49; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_50; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_51; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_52; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_53; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_54; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_55; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_56; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_57; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_58; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_59; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_60; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_61; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_62; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_63; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_64; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_65; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_66; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_67; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_68; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_69; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_70; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_71; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_72; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_73; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_74; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_75; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_76; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_77; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_78; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_79; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_80; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_81; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_82; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_83; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_84; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_85; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_86; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_87; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_88; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_89; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_90; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_91; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_92; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_93; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_94; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_95; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_96; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_97; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_98; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_99; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_100; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_101; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_102; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_103; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_104; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_105; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_106; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_107; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_108; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_109; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_110; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_111; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_112; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_113; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_114; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_115; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_116; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_117; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_118; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_119; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_120; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_121; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_122; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_123; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_124; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_125; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_126; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_127; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_128; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_129; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_130; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_131; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_132; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_133; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_134; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_135; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_136; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_137; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_138; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_139; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_140; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_141; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_142; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_143; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_144; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_145; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_146; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_147; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_148; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_149; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_150; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_151; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_152; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_153; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_154; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_155; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_156; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_157; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_158; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_159; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_160; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_161; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_162; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_163; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_164; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_165; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_166; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_167; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_168; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_169; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_170; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_171; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_172; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_173; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_174; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_175; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_176; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_177; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_178; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_179; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_180; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_181; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_182; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_183; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_184; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_185; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_186; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_187; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_188; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_189; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_190; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_191; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_192; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_193; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_194; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_195; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_196; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_197; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_198; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_199; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_200; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_201; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_202; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_203; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_204; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_205; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_206; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_207; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_208; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_209; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_210; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_211; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_212; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_213; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_214; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_215; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_216; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_217; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_218; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_219; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_220; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_221; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_222; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_223; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_224; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_225; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_226; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_227; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_228; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_229; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_230; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_231; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_232; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_233; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_234; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_235; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_236; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_237; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_238; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_239; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_240; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_241; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_242; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_243; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_244; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_245; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_246; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_247; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_248; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_249; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_250; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_251; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_252; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_253; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_254; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_255; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_256; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_257; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_258; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_259; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_260; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_261; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_262; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_263; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_264; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_265; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_266; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_267; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_268; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_269; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_270; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_271; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_272; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_273; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_274; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_275; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_276; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_277; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_278; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_279; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_280; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_281; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_282; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_283; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_284; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_285; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_286; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_287; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_288; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_289; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_290; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_291; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_292; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_293; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_294; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_295; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_296; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_297; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_298; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_299; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_300; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_301; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_302; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_303; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_304; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_305; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_306; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_307; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_308; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_309; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_310; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_311; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_312; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_313; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_314; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_315; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_316; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_317; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_318; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_319; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_320; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_321; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_322; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_323; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_324; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_325; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_326; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_327; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_328; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_329; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_330; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_331; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_332; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_333; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_334; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_335; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_336; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_337; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_338; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_339; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_340; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_341; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_342; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_343; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_344; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_345; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_346; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_347; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_348; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_349; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_350; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_351; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_352; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_353; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_354; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_355; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_356; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_357; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_358; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_359; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_360; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_361; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_362; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_363; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_364; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_365; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_366; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_367; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_368; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_369; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_370; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_371; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_372; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_373; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_374; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_375; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_376; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_377; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_378; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_379; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_380; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_381; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_382; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_383; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_384; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_385; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_386; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_387; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_388; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_389; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_390; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_391; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_392; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_393; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_394; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_395; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_396; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_397; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_398; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_399; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_400; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_401; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_402; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_403; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_404; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_405; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_406; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_407; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_408; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_409; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_410; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_411; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_412; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_413; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_414; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_415; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_416; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_417; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_418; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_419; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_420; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_421; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_422; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_423; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_424; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_425; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_426; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_427; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_428; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_429; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_430; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_431; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_432; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_433; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_434; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_435; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_436; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_437; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_438; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_439; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_440; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_441; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_442; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_443; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_444; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_445; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_446; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_447; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_448; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_449; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_450; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_451; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_452; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_453; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_454; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_455; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_456; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_457; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_458; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_459; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_460; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_461; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_462; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_463; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_464; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_465; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_466; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_467; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_468; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_469; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_470; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_471; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_472; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_473; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_474; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_475; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_476; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_477; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_478; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_479; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_480; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_481; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_482; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_483; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_484; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_485; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_486; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_487; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_488; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_489; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_490; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_491; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_492; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_493; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_494; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_495; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_496; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_497; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_498; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_499; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_500; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_501; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_502; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_503; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_504; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_505; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_506; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_507; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_508; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_509; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_510; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_511; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_512; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_513; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_514; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_515; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_516; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_517; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_518; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_519; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_520; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_521; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_522; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_523; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_524; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_525; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_526; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_527; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_528; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_529; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_530; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_531; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_532; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_533; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_534; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_535; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_536; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_537; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_538; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_539; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_540; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_541; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_542; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_543; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_544; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_545; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_546; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_547; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_548; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_549; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_550; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_551; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_552; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_553; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_554; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_555; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_556; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_557; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_558; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_559; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_560; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_561; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_562; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_563; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_564; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_565; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_566; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_567; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_568; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_569; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_570; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_571; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_572; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_573; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_574; // @[acccel_top.scala 166:22]
  wire [7:0] conv_io_weight_win_33_575; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_0; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_1; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_2; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_3; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_4; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_5; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_6; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_bias_data_7; // @[acccel_top.scala 166:22]
  wire  conv_io_bias_valid; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_0; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_1; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_2; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_3; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_4; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_5; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_6; // @[acccel_top.scala 166:22]
  wire [17:0] conv_io_conv_o_7; // @[acccel_top.scala 166:22]
  wire  acc_clock; // @[acccel_top.scala 182:21]
  wire  acc_reset; // @[acccel_top.scala 182:21]
  wire  acc_io_prev_data_zero; // @[acccel_top.scala 182:21]
  wire  acc_io_curr_data_zero; // @[acccel_top.scala 182:21]
  wire  acc_io_read_en; // @[acccel_top.scala 182:21]
  wire  acc_io_write_en; // @[acccel_top.scala 182:21]
  wire [11:0] acc_io_read_addr; // @[acccel_top.scala 182:21]
  wire [11:0] acc_io_write_addr; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_0; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_1; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_2; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_3; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_4; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_5; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_6; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_curr_data_7; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_0; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_1; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_2; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_3; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_4; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_5; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_6; // @[acccel_top.scala 182:21]
  wire [17:0] acc_io_acc_result_7; // @[acccel_top.scala 182:21]
  wire  quant_clock; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_0; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_1; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_2; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_3; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_4; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_5; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_6; // @[acccel_top.scala 195:23]
  wire [17:0] quant_io_acc_result_7; // @[acccel_top.scala 195:23]
  wire [15:0] quant_io_scale; // @[acccel_top.scala 195:23]
  wire [3:0] quant_io_shift; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_zero_point; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_0; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_1; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_2; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_3; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_4; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_5; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_6; // @[acccel_top.scala 195:23]
  wire [7:0] quant_io_quant_result_7; // @[acccel_top.scala 195:23]
  wire  pool_ctrl_clock; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_reset; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_io_pool_enable; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_zero_point; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_io_pool_finish; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_0; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_1; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_2; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_3; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_4; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_5; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_6; // @[acccel_top.scala 234:27]
  wire [7:0] pool_ctrl_io_pool_input_7; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_io_last_data_of_row; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_io_pool_outdata_valid; // @[acccel_top.scala 234:27]
  wire [11:0] pool_ctrl_io_ofm_write_addr; // @[acccel_top.scala 234:27]
  wire  pool_ctrl_io_ofm_en_write; // @[acccel_top.scala 234:27]
  wire [11:0] pool_ctrl_io_ofm_read_addr; // @[acccel_top.scala 234:27]
  wire [63:0] pool_ctrl_io_ofm_read_bundle; // @[acccel_top.scala 234:27]
  wire [9:0] pool_ctrl_io_row; // @[acccel_top.scala 234:27]
  wire [9:0] pool_ctrl_io_col; // @[acccel_top.scala 234:27]
  wire  pool_clock; // @[acccel_top.scala 249:22]
  wire  pool_reset; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_0; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_1; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_2; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_3; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_4; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_5; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_6; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_input_7; // @[acccel_top.scala 249:22]
  wire  pool_io_last_data_of_row; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_0; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_1; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_2; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_3; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_4; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_5; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_6; // @[acccel_top.scala 249:22]
  wire [7:0] pool_io_output_7; // @[acccel_top.scala 249:22]
  wire  pool_io_outdata_valid; // @[acccel_top.scala 249:22]
  wire  bn_add_clock; // @[acccel_top.scala 276:24]
  wire  bn_add_reset; // @[acccel_top.scala 276:24]
  wire [10:0] bn_add_io_ifm_read_addr; // @[acccel_top.scala 276:24]
  wire  bn_add_io_ifm_addr_read_sel; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_0; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_1; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_2; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_3; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_4; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_5; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_6; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_ifm_read_data_7; // @[acccel_top.scala 276:24]
  wire [11:0] bn_add_io_ofm_write_addr; // @[acccel_top.scala 276:24]
  wire  bn_add_io_ofm_en_write; // @[acccel_top.scala 276:24]
  wire [11:0] bn_add_io_ofm_read_addr; // @[acccel_top.scala 276:24]
  wire [63:0] bn_add_io_ofm_write_data; // @[acccel_top.scala 276:24]
  wire [63:0] bn_add_io_ofm_read_data; // @[acccel_top.scala 276:24]
  wire [9:0] bn_add_io_col; // @[acccel_top.scala 276:24]
  wire [9:0] bn_add_io_row; // @[acccel_top.scala 276:24]
  wire  bn_add_io_bottleneck_add_enable; // @[acccel_top.scala 276:24]
  wire  bn_add_io_bottleneck_add_finish; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_0; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_1; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_2; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_3; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_4; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_5; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_6; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in0_7; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_0; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_1; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_2; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_3; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_4; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_5; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_6; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_in1_7; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_0; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_1; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_2; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_3; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_4; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_5; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_6; // @[acccel_top.scala 276:24]
  wire [7:0] bn_add_io_bn_add_result_7; // @[acccel_top.scala 276:24]
  wire  ofm_clock; // @[acccel_top.scala 303:21]
  wire [11:0] ofm_io_bram_write_addr; // @[acccel_top.scala 303:21]
  wire  ofm_io_bram_en_write; // @[acccel_top.scala 303:21]
  wire [11:0] ofm_io_bram_read_addr; // @[acccel_top.scala 303:21]
  wire [63:0] ofm_io_ofm_store_bundle; // @[acccel_top.scala 303:21]
  wire [63:0] ofm_io_ofm_out_bundle; // @[acccel_top.scala 303:21]
  reg  bottleneck_work; // @[acccel_top.scala 88:34]
  reg  bottleneck_work_REG; // @[utils.scala 10:17]
  wire  _bottleneck_work_T_1 = ~bottleneck_work_REG & io_bottleneck_add_enable; // @[utils.scala 10:27]
  reg  bottleneck_work_REG_1; // @[utils.scala 10:17]
  wire  bottleneck_add_finish = bn_add_io_bottleneck_add_finish; // @[acccel_top.scala 279:27 89:37]
  wire  _bottleneck_work_T_3 = ~bottleneck_work_REG_1 & bottleneck_add_finish; // @[utils.scala 10:27]
  wire  _bottleneck_work_T_4 = _bottleneck_work_T_3 ? 1'h0 : bottleneck_work; // @[acccel_top.scala 90:75]
  wire [11:0] bn_add_ifm_read_addr = {{1'd0}, bn_add_io_ifm_read_addr}; // @[acccel_top.scala 286:26 91:36]
  wire [11:0] _ifm_buf_io_ifmbuf_bram_addr_read_s1_T = bottleneck_work ? bn_add_ifm_read_addr : {{1'd0},
    io_ifmbuf_bram_addr_read_s1}; // @[acccel_top.scala 96:47]
  wire  bn_add_ifm_addr_read_sel = bn_add_io_ifm_addr_read_sel; // @[acccel_top.scala 287:30 92:38]
  wire [31:0] ifmstream_0 = ifm_buf_io_ifm_o_data_0; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_0_lo = {sub_zero_io_data_out_1,sub_zero_io_data_out_0}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_0_hi = {sub_zero_io_data_out_3,sub_zero_io_data_out_2}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_1 = ifm_buf_io_ifm_o_data_1; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_1_lo = {sub_zero_io_data_out_5,sub_zero_io_data_out_4}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_1_hi = {sub_zero_io_data_out_7,sub_zero_io_data_out_6}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_2 = ifm_buf_io_ifm_o_data_2; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_2_lo = {sub_zero_io_data_out_9,sub_zero_io_data_out_8}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_2_hi = {sub_zero_io_data_out_11,sub_zero_io_data_out_10}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_3 = ifm_buf_io_ifm_o_data_3; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_3_lo = {sub_zero_io_data_out_13,sub_zero_io_data_out_12}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_3_hi = {sub_zero_io_data_out_15,sub_zero_io_data_out_14}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_4 = ifm_buf_io_ifm_o_data_4; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_4_lo = {sub_zero_io_data_out_17,sub_zero_io_data_out_16}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_4_hi = {sub_zero_io_data_out_19,sub_zero_io_data_out_18}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_5 = ifm_buf_io_ifm_o_data_5; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_5_lo = {sub_zero_io_data_out_21,sub_zero_io_data_out_20}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_5_hi = {sub_zero_io_data_out_23,sub_zero_io_data_out_22}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_6 = ifm_buf_io_ifm_o_data_6; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_6_lo = {sub_zero_io_data_out_25,sub_zero_io_data_out_24}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_6_hi = {sub_zero_io_data_out_27,sub_zero_io_data_out_26}; // @[Cat.scala 33:92]
  wire [31:0] ifmstream_7 = ifm_buf_io_ifm_o_data_7; // @[acccel_top.scala 116:22 94:25]
  wire [15:0] ifmstream_sub_zp_7_lo = {sub_zero_io_data_out_29,sub_zero_io_data_out_28}; // @[Cat.scala 33:92]
  wire [15:0] ifmstream_sub_zp_7_hi = {sub_zero_io_data_out_31,sub_zero_io_data_out_30}; // @[Cat.scala 33:92]
  wire [71:0] weight_win_0 = weight_buf_io_weight_out_0; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_1 = weight_buf_io_weight_out_1; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_2 = weight_buf_io_weight_out_2; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_3 = weight_buf_io_weight_out_3; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_4 = weight_buf_io_weight_out_4; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_5 = weight_buf_io_weight_out_5; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_6 = weight_buf_io_weight_out_6; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_7 = weight_buf_io_weight_out_7; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_8 = weight_buf_io_weight_out_8; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_9 = weight_buf_io_weight_out_9; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_10 = weight_buf_io_weight_out_10; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_11 = weight_buf_io_weight_out_11; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_12 = weight_buf_io_weight_out_12; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_13 = weight_buf_io_weight_out_13; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_14 = weight_buf_io_weight_out_14; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_15 = weight_buf_io_weight_out_15; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_16 = weight_buf_io_weight_out_16; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_17 = weight_buf_io_weight_out_17; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_18 = weight_buf_io_weight_out_18; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_19 = weight_buf_io_weight_out_19; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_20 = weight_buf_io_weight_out_20; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_21 = weight_buf_io_weight_out_21; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_22 = weight_buf_io_weight_out_22; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_23 = weight_buf_io_weight_out_23; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_24 = weight_buf_io_weight_out_24; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_25 = weight_buf_io_weight_out_25; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_26 = weight_buf_io_weight_out_26; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_27 = weight_buf_io_weight_out_27; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_28 = weight_buf_io_weight_out_28; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_29 = weight_buf_io_weight_out_29; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_30 = weight_buf_io_weight_out_30; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_31 = weight_buf_io_weight_out_31; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_32 = weight_buf_io_weight_out_32; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_33 = weight_buf_io_weight_out_33; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_34 = weight_buf_io_weight_out_34; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_35 = weight_buf_io_weight_out_35; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_36 = weight_buf_io_weight_out_36; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_37 = weight_buf_io_weight_out_37; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_38 = weight_buf_io_weight_out_38; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_39 = weight_buf_io_weight_out_39; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_40 = weight_buf_io_weight_out_40; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_41 = weight_buf_io_weight_out_41; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_42 = weight_buf_io_weight_out_42; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_43 = weight_buf_io_weight_out_43; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_44 = weight_buf_io_weight_out_44; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_45 = weight_buf_io_weight_out_45; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_46 = weight_buf_io_weight_out_46; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_47 = weight_buf_io_weight_out_47; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_48 = weight_buf_io_weight_out_48; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_49 = weight_buf_io_weight_out_49; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_50 = weight_buf_io_weight_out_50; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_51 = weight_buf_io_weight_out_51; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_52 = weight_buf_io_weight_out_52; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_53 = weight_buf_io_weight_out_53; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_54 = weight_buf_io_weight_out_54; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_55 = weight_buf_io_weight_out_55; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_56 = weight_buf_io_weight_out_56; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_57 = weight_buf_io_weight_out_57; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_58 = weight_buf_io_weight_out_58; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_59 = weight_buf_io_weight_out_59; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_60 = weight_buf_io_weight_out_60; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_61 = weight_buf_io_weight_out_61; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_62 = weight_buf_io_weight_out_62; // @[acccel_top.scala 119:26 129:38]
  wire [71:0] weight_win_63 = weight_buf_io_weight_out_63; // @[acccel_top.scala 119:26 129:38]
  wire [7:0] quant_result_0 = quant_io_quant_result_0; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_0 = io_skip_act ? quant_result_0 : io_act_outdata_0; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_1 = quant_io_quant_result_1; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_1 = io_skip_act ? quant_result_1 : io_act_outdata_1; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_2 = quant_io_quant_result_2; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_2 = io_skip_act ? quant_result_2 : io_act_outdata_2; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_3 = quant_io_quant_result_3; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_3 = io_skip_act ? quant_result_3 : io_act_outdata_3; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_4 = quant_io_quant_result_4; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_4 = io_skip_act ? quant_result_4 : io_act_outdata_4; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_5 = quant_io_quant_result_5; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_5 = io_skip_act ? quant_result_5 : io_act_outdata_5; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_6 = quant_io_quant_result_6; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_6 = io_skip_act ? quant_result_6 : io_act_outdata_6; // @[acccel_top.scala 257:24]
  wire [7:0] quant_result_7 = quant_io_quant_result_7; // @[acccel_top.scala 194:28 201:25]
  wire [7:0] conv_data_7 = io_skip_act ? quant_result_7 : io_act_outdata_7; // @[acccel_top.scala 257:24]
  wire [55:0] _ofm_conv_data_T_5 = {conv_data_6,conv_data_5,conv_data_4,conv_data_3,conv_data_2,conv_data_1,conv_data_0}
    ; // @[Cat.scala 33:92]
  wire [63:0] ofm_conv_data = {conv_data_7,conv_data_6,conv_data_5,conv_data_4,conv_data_3,conv_data_2,conv_data_1,
    conv_data_0}; // @[Cat.scala 33:92]
  wire [7:0] pool_output_1 = pool_io_output_1; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_0 = pool_io_output_0; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_2 = pool_io_output_2; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_3 = pool_io_output_3; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_4 = pool_io_output_4; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_5 = pool_io_output_5; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_6 = pool_io_output_6; // @[acccel_top.scala 230:27 254:24]
  wire [7:0] pool_output_7 = pool_io_output_7; // @[acccel_top.scala 230:27 254:24]
  wire [63:0] pool_data_bundle = {pool_output_7,pool_output_6,pool_output_5,pool_output_4,pool_output_3,pool_output_2,
    pool_output_1,pool_output_0}; // @[Cat.scala 33:92]
  reg  pool_work; // @[acccel_top.scala 294:28]
  reg  pool_work_REG; // @[utils.scala 10:17]
  wire  _pool_work_T_1 = ~pool_work_REG & io_pool_enable; // @[utils.scala 10:27]
  reg  pool_work_REG_1; // @[utils.scala 10:17]
  wire  pool_finish = pool_ctrl_io_pool_finish; // @[acccel_top.scala 231:25 237:17]
  wire  _pool_work_T_3 = ~pool_work_REG_1 & pool_finish; // @[utils.scala 10:27]
  wire  _pool_work_T_4 = _pool_work_T_3 ? 1'h0 : pool_work; // @[acccel_top.scala 295:59]
  wire [63:0] ofm_write_data = io_yolo_cls_en ? io_yolo_cls_data_after_compare : ofm_conv_data; // @[acccel_top.scala 297:27]
  wire [11:0] bn_add_ofm_write_addr = bn_add_io_ofm_write_addr; // @[acccel_top.scala 266:37 281:27]
  wire [11:0] _ofm_write_addr_T = bottleneck_work ? bn_add_ofm_write_addr : io_ofmbuf_bram_write_addr; // @[acccel_top.scala 298:63]
  wire [11:0] pool_ofm_write_addr = pool_ctrl_io_ofm_write_addr; // @[acccel_top.scala 224:35 238:25]
  wire  bn_add_ofm_en_write = bn_add_io_ofm_en_write; // @[acccel_top.scala 267:35 282:25]
  wire  _ofm_en_write_T = bottleneck_work ? bn_add_ofm_en_write : io_ofmbuf_bram_en_write; // @[acccel_top.scala 299:59]
  wire  pool_ofm_en_write = pool_ctrl_io_ofm_en_write; // @[acccel_top.scala 225:33 239:23]
  wire [11:0] bn_add_ofm_read_addr = bn_add_io_ofm_read_addr; // @[acccel_top.scala 268:36 283:26]
  wire [63:0] _ofm_read_addr_T = bottleneck_work ? {{52'd0}, bn_add_ofm_read_addr} : io_ofmbuf_bram_read_addr; // @[acccel_top.scala 300:61]
  wire [11:0] pool_ofm_read_addr = pool_ctrl_io_ofm_read_addr; // @[acccel_top.scala 227:34 241:24]
  wire [63:0] ofm_read_addr = pool_work ? {{52'd0}, pool_ofm_read_addr} : _ofm_read_addr_T; // @[acccel_top.scala 300:28]
  wire [63:0] bn_add_ofm_write_data = bn_add_io_ofm_write_data; // @[acccel_top.scala 269:37 284:27]
  wire [63:0] _ofm_store_bundle_T = bottleneck_work ? bn_add_ofm_write_data : ofm_write_data; // @[acccel_top.scala 301:64]
  IfmBuffer ifm_buf ( // @[acccel_top.scala 95:25]
    .clock(ifm_buf_clock),
    .reset(ifm_buf_reset),
    .io_ifmbuf_bram_addr_read_s1(ifm_buf_io_ifmbuf_bram_addr_read_s1),
    .io_ifmbuf_bram_addr_read_sel_s1(ifm_buf_io_ifmbuf_bram_addr_read_sel_s1),
    .io_ifmbuf_bram_addr_read_s2_singal(ifm_buf_io_ifmbuf_bram_addr_read_s2_singal),
    .io_ifmbuf_bram_addr_read_s2_double(ifm_buf_io_ifmbuf_bram_addr_read_s2_double),
    .io_bram_en_write(ifm_buf_io_bram_en_write),
    .io_upsample_enable(ifm_buf_io_upsample_enable),
    .io_recv_done(ifm_buf_io_recv_done),
    .io_buf_sel(ifm_buf_io_buf_sel),
    .io_s_mod(ifm_buf_io_s_mod),
    .io_col(ifm_buf_io_col),
    .io_in_0(ifm_buf_io_in_0),
    .io_in_1(ifm_buf_io_in_1),
    .io_in_2(ifm_buf_io_in_2),
    .io_in_3(ifm_buf_io_in_3),
    .io_in_4(ifm_buf_io_in_4),
    .io_in_5(ifm_buf_io_in_5),
    .io_in_6(ifm_buf_io_in_6),
    .io_in_7(ifm_buf_io_in_7),
    .io_ifm_o_data_0(ifm_buf_io_ifm_o_data_0),
    .io_ifm_o_data_1(ifm_buf_io_ifm_o_data_1),
    .io_ifm_o_data_2(ifm_buf_io_ifm_o_data_2),
    .io_ifm_o_data_3(ifm_buf_io_ifm_o_data_3),
    .io_ifm_o_data_4(ifm_buf_io_ifm_o_data_4),
    .io_ifm_o_data_5(ifm_buf_io_ifm_o_data_5),
    .io_ifm_o_data_6(ifm_buf_io_ifm_o_data_6),
    .io_ifm_o_data_7(ifm_buf_io_ifm_o_data_7),
    .io_pad_top(ifm_buf_io_pad_top),
    .io_pad_bottom(ifm_buf_io_pad_bottom),
    .io_pad_left_and_right(ifm_buf_io_pad_left_and_right),
    .io_zero_pad_valid_s2(ifm_buf_io_zero_pad_valid_s2),
    .io_zero_pad_valid_s1(ifm_buf_io_zero_pad_valid_s1),
    .io_zero_point_in(ifm_buf_io_zero_point_in)
  );
  WeightBuffer weight_buf ( // @[acccel_top.scala 120:28]
    .clock(weight_buf_clock),
    .reset(weight_buf_reset),
    .io_clear(weight_buf_io_clear),
    .io_bram_write_en(weight_buf_io_bram_write_en),
    .io_in_0(weight_buf_io_in_0),
    .io_in_1(weight_buf_io_in_1),
    .io_in_2(weight_buf_io_in_2),
    .io_in_3(weight_buf_io_in_3),
    .io_in_4(weight_buf_io_in_4),
    .io_in_5(weight_buf_io_in_5),
    .io_in_6(weight_buf_io_in_6),
    .io_in_7(weight_buf_io_in_7),
    .io_read_addr(weight_buf_io_read_addr),
    .io_sel_when_kernal_is_1(weight_buf_io_sel_when_kernal_is_1),
    .io_weight_out_0(weight_buf_io_weight_out_0),
    .io_weight_out_1(weight_buf_io_weight_out_1),
    .io_weight_out_2(weight_buf_io_weight_out_2),
    .io_weight_out_3(weight_buf_io_weight_out_3),
    .io_weight_out_4(weight_buf_io_weight_out_4),
    .io_weight_out_5(weight_buf_io_weight_out_5),
    .io_weight_out_6(weight_buf_io_weight_out_6),
    .io_weight_out_7(weight_buf_io_weight_out_7),
    .io_weight_out_8(weight_buf_io_weight_out_8),
    .io_weight_out_9(weight_buf_io_weight_out_9),
    .io_weight_out_10(weight_buf_io_weight_out_10),
    .io_weight_out_11(weight_buf_io_weight_out_11),
    .io_weight_out_12(weight_buf_io_weight_out_12),
    .io_weight_out_13(weight_buf_io_weight_out_13),
    .io_weight_out_14(weight_buf_io_weight_out_14),
    .io_weight_out_15(weight_buf_io_weight_out_15),
    .io_weight_out_16(weight_buf_io_weight_out_16),
    .io_weight_out_17(weight_buf_io_weight_out_17),
    .io_weight_out_18(weight_buf_io_weight_out_18),
    .io_weight_out_19(weight_buf_io_weight_out_19),
    .io_weight_out_20(weight_buf_io_weight_out_20),
    .io_weight_out_21(weight_buf_io_weight_out_21),
    .io_weight_out_22(weight_buf_io_weight_out_22),
    .io_weight_out_23(weight_buf_io_weight_out_23),
    .io_weight_out_24(weight_buf_io_weight_out_24),
    .io_weight_out_25(weight_buf_io_weight_out_25),
    .io_weight_out_26(weight_buf_io_weight_out_26),
    .io_weight_out_27(weight_buf_io_weight_out_27),
    .io_weight_out_28(weight_buf_io_weight_out_28),
    .io_weight_out_29(weight_buf_io_weight_out_29),
    .io_weight_out_30(weight_buf_io_weight_out_30),
    .io_weight_out_31(weight_buf_io_weight_out_31),
    .io_weight_out_32(weight_buf_io_weight_out_32),
    .io_weight_out_33(weight_buf_io_weight_out_33),
    .io_weight_out_34(weight_buf_io_weight_out_34),
    .io_weight_out_35(weight_buf_io_weight_out_35),
    .io_weight_out_36(weight_buf_io_weight_out_36),
    .io_weight_out_37(weight_buf_io_weight_out_37),
    .io_weight_out_38(weight_buf_io_weight_out_38),
    .io_weight_out_39(weight_buf_io_weight_out_39),
    .io_weight_out_40(weight_buf_io_weight_out_40),
    .io_weight_out_41(weight_buf_io_weight_out_41),
    .io_weight_out_42(weight_buf_io_weight_out_42),
    .io_weight_out_43(weight_buf_io_weight_out_43),
    .io_weight_out_44(weight_buf_io_weight_out_44),
    .io_weight_out_45(weight_buf_io_weight_out_45),
    .io_weight_out_46(weight_buf_io_weight_out_46),
    .io_weight_out_47(weight_buf_io_weight_out_47),
    .io_weight_out_48(weight_buf_io_weight_out_48),
    .io_weight_out_49(weight_buf_io_weight_out_49),
    .io_weight_out_50(weight_buf_io_weight_out_50),
    .io_weight_out_51(weight_buf_io_weight_out_51),
    .io_weight_out_52(weight_buf_io_weight_out_52),
    .io_weight_out_53(weight_buf_io_weight_out_53),
    .io_weight_out_54(weight_buf_io_weight_out_54),
    .io_weight_out_55(weight_buf_io_weight_out_55),
    .io_weight_out_56(weight_buf_io_weight_out_56),
    .io_weight_out_57(weight_buf_io_weight_out_57),
    .io_weight_out_58(weight_buf_io_weight_out_58),
    .io_weight_out_59(weight_buf_io_weight_out_59),
    .io_weight_out_60(weight_buf_io_weight_out_60),
    .io_weight_out_61(weight_buf_io_weight_out_61),
    .io_weight_out_62(weight_buf_io_weight_out_62),
    .io_weight_out_63(weight_buf_io_weight_out_63),
    .io_kernal(weight_buf_io_kernal)
  );
  BiasBuffer bias_buf ( // @[acccel_top.scala 134:26]
    .clock(bias_buf_clock),
    .reset(bias_buf_reset),
    .io_clear(bias_buf_io_clear),
    .io_bias_in(bias_buf_io_bias_in),
    .io_bram_addr_read(bias_buf_io_bram_addr_read),
    .io_bram_en_write(bias_buf_io_bram_en_write),
    .io_bias_data_0(bias_buf_io_bias_data_0),
    .io_bias_data_1(bias_buf_io_bias_data_1),
    .io_bias_data_2(bias_buf_io_bias_data_2),
    .io_bias_data_3(bias_buf_io_bias_data_3),
    .io_bias_data_4(bias_buf_io_bias_data_4),
    .io_bias_data_5(bias_buf_io_bias_data_5),
    .io_bias_data_6(bias_buf_io_bias_data_6),
    .io_bias_data_7(bias_buf_io_bias_data_7)
  );
  sub_zero_point sub_zero ( // @[acccel_top.scala 144:26]
    .clock(sub_zero_clock),
    .reset(sub_zero_reset),
    .io_zero_point(sub_zero_io_zero_point),
    .io_data_in_0(sub_zero_io_data_in_0),
    .io_data_in_1(sub_zero_io_data_in_1),
    .io_data_in_2(sub_zero_io_data_in_2),
    .io_data_in_3(sub_zero_io_data_in_3),
    .io_data_in_4(sub_zero_io_data_in_4),
    .io_data_in_5(sub_zero_io_data_in_5),
    .io_data_in_6(sub_zero_io_data_in_6),
    .io_data_in_7(sub_zero_io_data_in_7),
    .io_data_in_8(sub_zero_io_data_in_8),
    .io_data_in_9(sub_zero_io_data_in_9),
    .io_data_in_10(sub_zero_io_data_in_10),
    .io_data_in_11(sub_zero_io_data_in_11),
    .io_data_in_12(sub_zero_io_data_in_12),
    .io_data_in_13(sub_zero_io_data_in_13),
    .io_data_in_14(sub_zero_io_data_in_14),
    .io_data_in_15(sub_zero_io_data_in_15),
    .io_data_in_16(sub_zero_io_data_in_16),
    .io_data_in_17(sub_zero_io_data_in_17),
    .io_data_in_18(sub_zero_io_data_in_18),
    .io_data_in_19(sub_zero_io_data_in_19),
    .io_data_in_20(sub_zero_io_data_in_20),
    .io_data_in_21(sub_zero_io_data_in_21),
    .io_data_in_22(sub_zero_io_data_in_22),
    .io_data_in_23(sub_zero_io_data_in_23),
    .io_data_in_24(sub_zero_io_data_in_24),
    .io_data_in_25(sub_zero_io_data_in_25),
    .io_data_in_26(sub_zero_io_data_in_26),
    .io_data_in_27(sub_zero_io_data_in_27),
    .io_data_in_28(sub_zero_io_data_in_28),
    .io_data_in_29(sub_zero_io_data_in_29),
    .io_data_in_30(sub_zero_io_data_in_30),
    .io_data_in_31(sub_zero_io_data_in_31),
    .io_data_out_0(sub_zero_io_data_out_0),
    .io_data_out_1(sub_zero_io_data_out_1),
    .io_data_out_2(sub_zero_io_data_out_2),
    .io_data_out_3(sub_zero_io_data_out_3),
    .io_data_out_4(sub_zero_io_data_out_4),
    .io_data_out_5(sub_zero_io_data_out_5),
    .io_data_out_6(sub_zero_io_data_out_6),
    .io_data_out_7(sub_zero_io_data_out_7),
    .io_data_out_8(sub_zero_io_data_out_8),
    .io_data_out_9(sub_zero_io_data_out_9),
    .io_data_out_10(sub_zero_io_data_out_10),
    .io_data_out_11(sub_zero_io_data_out_11),
    .io_data_out_12(sub_zero_io_data_out_12),
    .io_data_out_13(sub_zero_io_data_out_13),
    .io_data_out_14(sub_zero_io_data_out_14),
    .io_data_out_15(sub_zero_io_data_out_15),
    .io_data_out_16(sub_zero_io_data_out_16),
    .io_data_out_17(sub_zero_io_data_out_17),
    .io_data_out_18(sub_zero_io_data_out_18),
    .io_data_out_19(sub_zero_io_data_out_19),
    .io_data_out_20(sub_zero_io_data_out_20),
    .io_data_out_21(sub_zero_io_data_out_21),
    .io_data_out_22(sub_zero_io_data_out_22),
    .io_data_out_23(sub_zero_io_data_out_23),
    .io_data_out_24(sub_zero_io_data_out_24),
    .io_data_out_25(sub_zero_io_data_out_25),
    .io_data_out_26(sub_zero_io_data_out_26),
    .io_data_out_27(sub_zero_io_data_out_27),
    .io_data_out_28(sub_zero_io_data_out_28),
    .io_data_out_29(sub_zero_io_data_out_29),
    .io_data_out_30(sub_zero_io_data_out_30),
    .io_data_out_31(sub_zero_io_data_out_31)
  );
  LineBuffer_extend line_buf ( // @[acccel_top.scala 154:26]
    .clock(line_buf_clock),
    .reset(line_buf_reset),
    .io_sel(line_buf_io_sel),
    .io_s_mod(line_buf_io_s_mod),
    .io_lineBuffer_i_data_0(line_buf_io_lineBuffer_i_data_0),
    .io_lineBuffer_i_data_1(line_buf_io_lineBuffer_i_data_1),
    .io_lineBuffer_i_data_2(line_buf_io_lineBuffer_i_data_2),
    .io_lineBuffer_i_data_3(line_buf_io_lineBuffer_i_data_3),
    .io_lineBuffer_i_data_4(line_buf_io_lineBuffer_i_data_4),
    .io_lineBuffer_i_data_5(line_buf_io_lineBuffer_i_data_5),
    .io_lineBuffer_i_data_6(line_buf_io_lineBuffer_i_data_6),
    .io_lineBuffer_i_data_7(line_buf_io_lineBuffer_i_data_7),
    .io_lineBuffer_o_data_0(line_buf_io_lineBuffer_o_data_0),
    .io_lineBuffer_o_data_1(line_buf_io_lineBuffer_o_data_1),
    .io_lineBuffer_o_data_2(line_buf_io_lineBuffer_o_data_2),
    .io_lineBuffer_o_data_3(line_buf_io_lineBuffer_o_data_3),
    .io_lineBuffer_o_data_4(line_buf_io_lineBuffer_o_data_4),
    .io_lineBuffer_o_data_5(line_buf_io_lineBuffer_o_data_5),
    .io_lineBuffer_o_data_6(line_buf_io_lineBuffer_o_data_6),
    .io_lineBuffer_o_data_7(line_buf_io_lineBuffer_o_data_7),
    .io_lineBuffer_o_data_8(line_buf_io_lineBuffer_o_data_8),
    .io_lineBuffer_o_data_9(line_buf_io_lineBuffer_o_data_9),
    .io_lineBuffer_o_data_10(line_buf_io_lineBuffer_o_data_10),
    .io_lineBuffer_o_data_11(line_buf_io_lineBuffer_o_data_11),
    .io_lineBuffer_o_data_12(line_buf_io_lineBuffer_o_data_12),
    .io_lineBuffer_o_data_13(line_buf_io_lineBuffer_o_data_13),
    .io_lineBuffer_o_data_14(line_buf_io_lineBuffer_o_data_14),
    .io_lineBuffer_o_data_15(line_buf_io_lineBuffer_o_data_15),
    .io_lineBuffer_o_data_16(line_buf_io_lineBuffer_o_data_16),
    .io_lineBuffer_o_data_17(line_buf_io_lineBuffer_o_data_17),
    .io_lineBuffer_o_data_18(line_buf_io_lineBuffer_o_data_18),
    .io_lineBuffer_o_data_19(line_buf_io_lineBuffer_o_data_19),
    .io_lineBuffer_o_data_20(line_buf_io_lineBuffer_o_data_20),
    .io_lineBuffer_o_data_21(line_buf_io_lineBuffer_o_data_21),
    .io_lineBuffer_o_data_22(line_buf_io_lineBuffer_o_data_22),
    .io_lineBuffer_o_data_23(line_buf_io_lineBuffer_o_data_23),
    .io_lineBuffer_o_data_24(line_buf_io_lineBuffer_o_data_24),
    .io_lineBuffer_o_data_25(line_buf_io_lineBuffer_o_data_25),
    .io_lineBuffer_o_data_26(line_buf_io_lineBuffer_o_data_26),
    .io_lineBuffer_o_data_27(line_buf_io_lineBuffer_o_data_27),
    .io_lineBuffer_o_data_28(line_buf_io_lineBuffer_o_data_28),
    .io_lineBuffer_o_data_29(line_buf_io_lineBuffer_o_data_29),
    .io_lineBuffer_o_data_30(line_buf_io_lineBuffer_o_data_30),
    .io_lineBuffer_o_data_31(line_buf_io_lineBuffer_o_data_31),
    .io_lineBuffer_o_data_32(line_buf_io_lineBuffer_o_data_32),
    .io_lineBuffer_o_data_33(line_buf_io_lineBuffer_o_data_33),
    .io_lineBuffer_o_data_34(line_buf_io_lineBuffer_o_data_34),
    .io_lineBuffer_o_data_35(line_buf_io_lineBuffer_o_data_35),
    .io_lineBuffer_o_data_36(line_buf_io_lineBuffer_o_data_36),
    .io_lineBuffer_o_data_37(line_buf_io_lineBuffer_o_data_37),
    .io_lineBuffer_o_data_38(line_buf_io_lineBuffer_o_data_38),
    .io_lineBuffer_o_data_39(line_buf_io_lineBuffer_o_data_39),
    .io_lineBuffer_o_data_40(line_buf_io_lineBuffer_o_data_40),
    .io_lineBuffer_o_data_41(line_buf_io_lineBuffer_o_data_41),
    .io_lineBuffer_o_data_42(line_buf_io_lineBuffer_o_data_42),
    .io_lineBuffer_o_data_43(line_buf_io_lineBuffer_o_data_43),
    .io_lineBuffer_o_data_44(line_buf_io_lineBuffer_o_data_44),
    .io_lineBuffer_o_data_45(line_buf_io_lineBuffer_o_data_45),
    .io_lineBuffer_o_data_46(line_buf_io_lineBuffer_o_data_46),
    .io_lineBuffer_o_data_47(line_buf_io_lineBuffer_o_data_47),
    .io_lineBuffer_o_data_48(line_buf_io_lineBuffer_o_data_48),
    .io_lineBuffer_o_data_49(line_buf_io_lineBuffer_o_data_49),
    .io_lineBuffer_o_data_50(line_buf_io_lineBuffer_o_data_50),
    .io_lineBuffer_o_data_51(line_buf_io_lineBuffer_o_data_51),
    .io_lineBuffer_o_data_52(line_buf_io_lineBuffer_o_data_52),
    .io_lineBuffer_o_data_53(line_buf_io_lineBuffer_o_data_53),
    .io_lineBuffer_o_data_54(line_buf_io_lineBuffer_o_data_54),
    .io_lineBuffer_o_data_55(line_buf_io_lineBuffer_o_data_55),
    .io_lineBuffer_o_data_56(line_buf_io_lineBuffer_o_data_56),
    .io_lineBuffer_o_data_57(line_buf_io_lineBuffer_o_data_57),
    .io_lineBuffer_o_data_58(line_buf_io_lineBuffer_o_data_58),
    .io_lineBuffer_o_data_59(line_buf_io_lineBuffer_o_data_59),
    .io_lineBuffer_o_data_60(line_buf_io_lineBuffer_o_data_60),
    .io_lineBuffer_o_data_61(line_buf_io_lineBuffer_o_data_61),
    .io_lineBuffer_o_data_62(line_buf_io_lineBuffer_o_data_62),
    .io_lineBuffer_o_data_63(line_buf_io_lineBuffer_o_data_63),
    .io_lineBuffer_o_data_64(line_buf_io_lineBuffer_o_data_64),
    .io_lineBuffer_o_data_65(line_buf_io_lineBuffer_o_data_65),
    .io_lineBuffer_o_data_66(line_buf_io_lineBuffer_o_data_66),
    .io_lineBuffer_o_data_67(line_buf_io_lineBuffer_o_data_67),
    .io_lineBuffer_o_data_68(line_buf_io_lineBuffer_o_data_68),
    .io_lineBuffer_o_data_69(line_buf_io_lineBuffer_o_data_69),
    .io_lineBuffer_o_data_70(line_buf_io_lineBuffer_o_data_70),
    .io_lineBuffer_o_data_71(line_buf_io_lineBuffer_o_data_71)
  );
  Conv conv ( // @[acccel_top.scala 166:22]
    .clock(conv_clock),
    .io_ifm_win_33_0(conv_io_ifm_win_33_0),
    .io_ifm_win_33_1(conv_io_ifm_win_33_1),
    .io_ifm_win_33_2(conv_io_ifm_win_33_2),
    .io_ifm_win_33_3(conv_io_ifm_win_33_3),
    .io_ifm_win_33_4(conv_io_ifm_win_33_4),
    .io_ifm_win_33_5(conv_io_ifm_win_33_5),
    .io_ifm_win_33_6(conv_io_ifm_win_33_6),
    .io_ifm_win_33_7(conv_io_ifm_win_33_7),
    .io_ifm_win_33_8(conv_io_ifm_win_33_8),
    .io_ifm_win_33_9(conv_io_ifm_win_33_9),
    .io_ifm_win_33_10(conv_io_ifm_win_33_10),
    .io_ifm_win_33_11(conv_io_ifm_win_33_11),
    .io_ifm_win_33_12(conv_io_ifm_win_33_12),
    .io_ifm_win_33_13(conv_io_ifm_win_33_13),
    .io_ifm_win_33_14(conv_io_ifm_win_33_14),
    .io_ifm_win_33_15(conv_io_ifm_win_33_15),
    .io_ifm_win_33_16(conv_io_ifm_win_33_16),
    .io_ifm_win_33_17(conv_io_ifm_win_33_17),
    .io_ifm_win_33_18(conv_io_ifm_win_33_18),
    .io_ifm_win_33_19(conv_io_ifm_win_33_19),
    .io_ifm_win_33_20(conv_io_ifm_win_33_20),
    .io_ifm_win_33_21(conv_io_ifm_win_33_21),
    .io_ifm_win_33_22(conv_io_ifm_win_33_22),
    .io_ifm_win_33_23(conv_io_ifm_win_33_23),
    .io_ifm_win_33_24(conv_io_ifm_win_33_24),
    .io_ifm_win_33_25(conv_io_ifm_win_33_25),
    .io_ifm_win_33_26(conv_io_ifm_win_33_26),
    .io_ifm_win_33_27(conv_io_ifm_win_33_27),
    .io_ifm_win_33_28(conv_io_ifm_win_33_28),
    .io_ifm_win_33_29(conv_io_ifm_win_33_29),
    .io_ifm_win_33_30(conv_io_ifm_win_33_30),
    .io_ifm_win_33_31(conv_io_ifm_win_33_31),
    .io_ifm_win_33_32(conv_io_ifm_win_33_32),
    .io_ifm_win_33_33(conv_io_ifm_win_33_33),
    .io_ifm_win_33_34(conv_io_ifm_win_33_34),
    .io_ifm_win_33_35(conv_io_ifm_win_33_35),
    .io_ifm_win_33_36(conv_io_ifm_win_33_36),
    .io_ifm_win_33_37(conv_io_ifm_win_33_37),
    .io_ifm_win_33_38(conv_io_ifm_win_33_38),
    .io_ifm_win_33_39(conv_io_ifm_win_33_39),
    .io_ifm_win_33_40(conv_io_ifm_win_33_40),
    .io_ifm_win_33_41(conv_io_ifm_win_33_41),
    .io_ifm_win_33_42(conv_io_ifm_win_33_42),
    .io_ifm_win_33_43(conv_io_ifm_win_33_43),
    .io_ifm_win_33_44(conv_io_ifm_win_33_44),
    .io_ifm_win_33_45(conv_io_ifm_win_33_45),
    .io_ifm_win_33_46(conv_io_ifm_win_33_46),
    .io_ifm_win_33_47(conv_io_ifm_win_33_47),
    .io_ifm_win_33_48(conv_io_ifm_win_33_48),
    .io_ifm_win_33_49(conv_io_ifm_win_33_49),
    .io_ifm_win_33_50(conv_io_ifm_win_33_50),
    .io_ifm_win_33_51(conv_io_ifm_win_33_51),
    .io_ifm_win_33_52(conv_io_ifm_win_33_52),
    .io_ifm_win_33_53(conv_io_ifm_win_33_53),
    .io_ifm_win_33_54(conv_io_ifm_win_33_54),
    .io_ifm_win_33_55(conv_io_ifm_win_33_55),
    .io_ifm_win_33_56(conv_io_ifm_win_33_56),
    .io_ifm_win_33_57(conv_io_ifm_win_33_57),
    .io_ifm_win_33_58(conv_io_ifm_win_33_58),
    .io_ifm_win_33_59(conv_io_ifm_win_33_59),
    .io_ifm_win_33_60(conv_io_ifm_win_33_60),
    .io_ifm_win_33_61(conv_io_ifm_win_33_61),
    .io_ifm_win_33_62(conv_io_ifm_win_33_62),
    .io_ifm_win_33_63(conv_io_ifm_win_33_63),
    .io_ifm_win_33_64(conv_io_ifm_win_33_64),
    .io_ifm_win_33_65(conv_io_ifm_win_33_65),
    .io_ifm_win_33_66(conv_io_ifm_win_33_66),
    .io_ifm_win_33_67(conv_io_ifm_win_33_67),
    .io_ifm_win_33_68(conv_io_ifm_win_33_68),
    .io_ifm_win_33_69(conv_io_ifm_win_33_69),
    .io_ifm_win_33_70(conv_io_ifm_win_33_70),
    .io_ifm_win_33_71(conv_io_ifm_win_33_71),
    .io_weight_win_33_0(conv_io_weight_win_33_0),
    .io_weight_win_33_1(conv_io_weight_win_33_1),
    .io_weight_win_33_2(conv_io_weight_win_33_2),
    .io_weight_win_33_3(conv_io_weight_win_33_3),
    .io_weight_win_33_4(conv_io_weight_win_33_4),
    .io_weight_win_33_5(conv_io_weight_win_33_5),
    .io_weight_win_33_6(conv_io_weight_win_33_6),
    .io_weight_win_33_7(conv_io_weight_win_33_7),
    .io_weight_win_33_8(conv_io_weight_win_33_8),
    .io_weight_win_33_9(conv_io_weight_win_33_9),
    .io_weight_win_33_10(conv_io_weight_win_33_10),
    .io_weight_win_33_11(conv_io_weight_win_33_11),
    .io_weight_win_33_12(conv_io_weight_win_33_12),
    .io_weight_win_33_13(conv_io_weight_win_33_13),
    .io_weight_win_33_14(conv_io_weight_win_33_14),
    .io_weight_win_33_15(conv_io_weight_win_33_15),
    .io_weight_win_33_16(conv_io_weight_win_33_16),
    .io_weight_win_33_17(conv_io_weight_win_33_17),
    .io_weight_win_33_18(conv_io_weight_win_33_18),
    .io_weight_win_33_19(conv_io_weight_win_33_19),
    .io_weight_win_33_20(conv_io_weight_win_33_20),
    .io_weight_win_33_21(conv_io_weight_win_33_21),
    .io_weight_win_33_22(conv_io_weight_win_33_22),
    .io_weight_win_33_23(conv_io_weight_win_33_23),
    .io_weight_win_33_24(conv_io_weight_win_33_24),
    .io_weight_win_33_25(conv_io_weight_win_33_25),
    .io_weight_win_33_26(conv_io_weight_win_33_26),
    .io_weight_win_33_27(conv_io_weight_win_33_27),
    .io_weight_win_33_28(conv_io_weight_win_33_28),
    .io_weight_win_33_29(conv_io_weight_win_33_29),
    .io_weight_win_33_30(conv_io_weight_win_33_30),
    .io_weight_win_33_31(conv_io_weight_win_33_31),
    .io_weight_win_33_32(conv_io_weight_win_33_32),
    .io_weight_win_33_33(conv_io_weight_win_33_33),
    .io_weight_win_33_34(conv_io_weight_win_33_34),
    .io_weight_win_33_35(conv_io_weight_win_33_35),
    .io_weight_win_33_36(conv_io_weight_win_33_36),
    .io_weight_win_33_37(conv_io_weight_win_33_37),
    .io_weight_win_33_38(conv_io_weight_win_33_38),
    .io_weight_win_33_39(conv_io_weight_win_33_39),
    .io_weight_win_33_40(conv_io_weight_win_33_40),
    .io_weight_win_33_41(conv_io_weight_win_33_41),
    .io_weight_win_33_42(conv_io_weight_win_33_42),
    .io_weight_win_33_43(conv_io_weight_win_33_43),
    .io_weight_win_33_44(conv_io_weight_win_33_44),
    .io_weight_win_33_45(conv_io_weight_win_33_45),
    .io_weight_win_33_46(conv_io_weight_win_33_46),
    .io_weight_win_33_47(conv_io_weight_win_33_47),
    .io_weight_win_33_48(conv_io_weight_win_33_48),
    .io_weight_win_33_49(conv_io_weight_win_33_49),
    .io_weight_win_33_50(conv_io_weight_win_33_50),
    .io_weight_win_33_51(conv_io_weight_win_33_51),
    .io_weight_win_33_52(conv_io_weight_win_33_52),
    .io_weight_win_33_53(conv_io_weight_win_33_53),
    .io_weight_win_33_54(conv_io_weight_win_33_54),
    .io_weight_win_33_55(conv_io_weight_win_33_55),
    .io_weight_win_33_56(conv_io_weight_win_33_56),
    .io_weight_win_33_57(conv_io_weight_win_33_57),
    .io_weight_win_33_58(conv_io_weight_win_33_58),
    .io_weight_win_33_59(conv_io_weight_win_33_59),
    .io_weight_win_33_60(conv_io_weight_win_33_60),
    .io_weight_win_33_61(conv_io_weight_win_33_61),
    .io_weight_win_33_62(conv_io_weight_win_33_62),
    .io_weight_win_33_63(conv_io_weight_win_33_63),
    .io_weight_win_33_64(conv_io_weight_win_33_64),
    .io_weight_win_33_65(conv_io_weight_win_33_65),
    .io_weight_win_33_66(conv_io_weight_win_33_66),
    .io_weight_win_33_67(conv_io_weight_win_33_67),
    .io_weight_win_33_68(conv_io_weight_win_33_68),
    .io_weight_win_33_69(conv_io_weight_win_33_69),
    .io_weight_win_33_70(conv_io_weight_win_33_70),
    .io_weight_win_33_71(conv_io_weight_win_33_71),
    .io_weight_win_33_72(conv_io_weight_win_33_72),
    .io_weight_win_33_73(conv_io_weight_win_33_73),
    .io_weight_win_33_74(conv_io_weight_win_33_74),
    .io_weight_win_33_75(conv_io_weight_win_33_75),
    .io_weight_win_33_76(conv_io_weight_win_33_76),
    .io_weight_win_33_77(conv_io_weight_win_33_77),
    .io_weight_win_33_78(conv_io_weight_win_33_78),
    .io_weight_win_33_79(conv_io_weight_win_33_79),
    .io_weight_win_33_80(conv_io_weight_win_33_80),
    .io_weight_win_33_81(conv_io_weight_win_33_81),
    .io_weight_win_33_82(conv_io_weight_win_33_82),
    .io_weight_win_33_83(conv_io_weight_win_33_83),
    .io_weight_win_33_84(conv_io_weight_win_33_84),
    .io_weight_win_33_85(conv_io_weight_win_33_85),
    .io_weight_win_33_86(conv_io_weight_win_33_86),
    .io_weight_win_33_87(conv_io_weight_win_33_87),
    .io_weight_win_33_88(conv_io_weight_win_33_88),
    .io_weight_win_33_89(conv_io_weight_win_33_89),
    .io_weight_win_33_90(conv_io_weight_win_33_90),
    .io_weight_win_33_91(conv_io_weight_win_33_91),
    .io_weight_win_33_92(conv_io_weight_win_33_92),
    .io_weight_win_33_93(conv_io_weight_win_33_93),
    .io_weight_win_33_94(conv_io_weight_win_33_94),
    .io_weight_win_33_95(conv_io_weight_win_33_95),
    .io_weight_win_33_96(conv_io_weight_win_33_96),
    .io_weight_win_33_97(conv_io_weight_win_33_97),
    .io_weight_win_33_98(conv_io_weight_win_33_98),
    .io_weight_win_33_99(conv_io_weight_win_33_99),
    .io_weight_win_33_100(conv_io_weight_win_33_100),
    .io_weight_win_33_101(conv_io_weight_win_33_101),
    .io_weight_win_33_102(conv_io_weight_win_33_102),
    .io_weight_win_33_103(conv_io_weight_win_33_103),
    .io_weight_win_33_104(conv_io_weight_win_33_104),
    .io_weight_win_33_105(conv_io_weight_win_33_105),
    .io_weight_win_33_106(conv_io_weight_win_33_106),
    .io_weight_win_33_107(conv_io_weight_win_33_107),
    .io_weight_win_33_108(conv_io_weight_win_33_108),
    .io_weight_win_33_109(conv_io_weight_win_33_109),
    .io_weight_win_33_110(conv_io_weight_win_33_110),
    .io_weight_win_33_111(conv_io_weight_win_33_111),
    .io_weight_win_33_112(conv_io_weight_win_33_112),
    .io_weight_win_33_113(conv_io_weight_win_33_113),
    .io_weight_win_33_114(conv_io_weight_win_33_114),
    .io_weight_win_33_115(conv_io_weight_win_33_115),
    .io_weight_win_33_116(conv_io_weight_win_33_116),
    .io_weight_win_33_117(conv_io_weight_win_33_117),
    .io_weight_win_33_118(conv_io_weight_win_33_118),
    .io_weight_win_33_119(conv_io_weight_win_33_119),
    .io_weight_win_33_120(conv_io_weight_win_33_120),
    .io_weight_win_33_121(conv_io_weight_win_33_121),
    .io_weight_win_33_122(conv_io_weight_win_33_122),
    .io_weight_win_33_123(conv_io_weight_win_33_123),
    .io_weight_win_33_124(conv_io_weight_win_33_124),
    .io_weight_win_33_125(conv_io_weight_win_33_125),
    .io_weight_win_33_126(conv_io_weight_win_33_126),
    .io_weight_win_33_127(conv_io_weight_win_33_127),
    .io_weight_win_33_128(conv_io_weight_win_33_128),
    .io_weight_win_33_129(conv_io_weight_win_33_129),
    .io_weight_win_33_130(conv_io_weight_win_33_130),
    .io_weight_win_33_131(conv_io_weight_win_33_131),
    .io_weight_win_33_132(conv_io_weight_win_33_132),
    .io_weight_win_33_133(conv_io_weight_win_33_133),
    .io_weight_win_33_134(conv_io_weight_win_33_134),
    .io_weight_win_33_135(conv_io_weight_win_33_135),
    .io_weight_win_33_136(conv_io_weight_win_33_136),
    .io_weight_win_33_137(conv_io_weight_win_33_137),
    .io_weight_win_33_138(conv_io_weight_win_33_138),
    .io_weight_win_33_139(conv_io_weight_win_33_139),
    .io_weight_win_33_140(conv_io_weight_win_33_140),
    .io_weight_win_33_141(conv_io_weight_win_33_141),
    .io_weight_win_33_142(conv_io_weight_win_33_142),
    .io_weight_win_33_143(conv_io_weight_win_33_143),
    .io_weight_win_33_144(conv_io_weight_win_33_144),
    .io_weight_win_33_145(conv_io_weight_win_33_145),
    .io_weight_win_33_146(conv_io_weight_win_33_146),
    .io_weight_win_33_147(conv_io_weight_win_33_147),
    .io_weight_win_33_148(conv_io_weight_win_33_148),
    .io_weight_win_33_149(conv_io_weight_win_33_149),
    .io_weight_win_33_150(conv_io_weight_win_33_150),
    .io_weight_win_33_151(conv_io_weight_win_33_151),
    .io_weight_win_33_152(conv_io_weight_win_33_152),
    .io_weight_win_33_153(conv_io_weight_win_33_153),
    .io_weight_win_33_154(conv_io_weight_win_33_154),
    .io_weight_win_33_155(conv_io_weight_win_33_155),
    .io_weight_win_33_156(conv_io_weight_win_33_156),
    .io_weight_win_33_157(conv_io_weight_win_33_157),
    .io_weight_win_33_158(conv_io_weight_win_33_158),
    .io_weight_win_33_159(conv_io_weight_win_33_159),
    .io_weight_win_33_160(conv_io_weight_win_33_160),
    .io_weight_win_33_161(conv_io_weight_win_33_161),
    .io_weight_win_33_162(conv_io_weight_win_33_162),
    .io_weight_win_33_163(conv_io_weight_win_33_163),
    .io_weight_win_33_164(conv_io_weight_win_33_164),
    .io_weight_win_33_165(conv_io_weight_win_33_165),
    .io_weight_win_33_166(conv_io_weight_win_33_166),
    .io_weight_win_33_167(conv_io_weight_win_33_167),
    .io_weight_win_33_168(conv_io_weight_win_33_168),
    .io_weight_win_33_169(conv_io_weight_win_33_169),
    .io_weight_win_33_170(conv_io_weight_win_33_170),
    .io_weight_win_33_171(conv_io_weight_win_33_171),
    .io_weight_win_33_172(conv_io_weight_win_33_172),
    .io_weight_win_33_173(conv_io_weight_win_33_173),
    .io_weight_win_33_174(conv_io_weight_win_33_174),
    .io_weight_win_33_175(conv_io_weight_win_33_175),
    .io_weight_win_33_176(conv_io_weight_win_33_176),
    .io_weight_win_33_177(conv_io_weight_win_33_177),
    .io_weight_win_33_178(conv_io_weight_win_33_178),
    .io_weight_win_33_179(conv_io_weight_win_33_179),
    .io_weight_win_33_180(conv_io_weight_win_33_180),
    .io_weight_win_33_181(conv_io_weight_win_33_181),
    .io_weight_win_33_182(conv_io_weight_win_33_182),
    .io_weight_win_33_183(conv_io_weight_win_33_183),
    .io_weight_win_33_184(conv_io_weight_win_33_184),
    .io_weight_win_33_185(conv_io_weight_win_33_185),
    .io_weight_win_33_186(conv_io_weight_win_33_186),
    .io_weight_win_33_187(conv_io_weight_win_33_187),
    .io_weight_win_33_188(conv_io_weight_win_33_188),
    .io_weight_win_33_189(conv_io_weight_win_33_189),
    .io_weight_win_33_190(conv_io_weight_win_33_190),
    .io_weight_win_33_191(conv_io_weight_win_33_191),
    .io_weight_win_33_192(conv_io_weight_win_33_192),
    .io_weight_win_33_193(conv_io_weight_win_33_193),
    .io_weight_win_33_194(conv_io_weight_win_33_194),
    .io_weight_win_33_195(conv_io_weight_win_33_195),
    .io_weight_win_33_196(conv_io_weight_win_33_196),
    .io_weight_win_33_197(conv_io_weight_win_33_197),
    .io_weight_win_33_198(conv_io_weight_win_33_198),
    .io_weight_win_33_199(conv_io_weight_win_33_199),
    .io_weight_win_33_200(conv_io_weight_win_33_200),
    .io_weight_win_33_201(conv_io_weight_win_33_201),
    .io_weight_win_33_202(conv_io_weight_win_33_202),
    .io_weight_win_33_203(conv_io_weight_win_33_203),
    .io_weight_win_33_204(conv_io_weight_win_33_204),
    .io_weight_win_33_205(conv_io_weight_win_33_205),
    .io_weight_win_33_206(conv_io_weight_win_33_206),
    .io_weight_win_33_207(conv_io_weight_win_33_207),
    .io_weight_win_33_208(conv_io_weight_win_33_208),
    .io_weight_win_33_209(conv_io_weight_win_33_209),
    .io_weight_win_33_210(conv_io_weight_win_33_210),
    .io_weight_win_33_211(conv_io_weight_win_33_211),
    .io_weight_win_33_212(conv_io_weight_win_33_212),
    .io_weight_win_33_213(conv_io_weight_win_33_213),
    .io_weight_win_33_214(conv_io_weight_win_33_214),
    .io_weight_win_33_215(conv_io_weight_win_33_215),
    .io_weight_win_33_216(conv_io_weight_win_33_216),
    .io_weight_win_33_217(conv_io_weight_win_33_217),
    .io_weight_win_33_218(conv_io_weight_win_33_218),
    .io_weight_win_33_219(conv_io_weight_win_33_219),
    .io_weight_win_33_220(conv_io_weight_win_33_220),
    .io_weight_win_33_221(conv_io_weight_win_33_221),
    .io_weight_win_33_222(conv_io_weight_win_33_222),
    .io_weight_win_33_223(conv_io_weight_win_33_223),
    .io_weight_win_33_224(conv_io_weight_win_33_224),
    .io_weight_win_33_225(conv_io_weight_win_33_225),
    .io_weight_win_33_226(conv_io_weight_win_33_226),
    .io_weight_win_33_227(conv_io_weight_win_33_227),
    .io_weight_win_33_228(conv_io_weight_win_33_228),
    .io_weight_win_33_229(conv_io_weight_win_33_229),
    .io_weight_win_33_230(conv_io_weight_win_33_230),
    .io_weight_win_33_231(conv_io_weight_win_33_231),
    .io_weight_win_33_232(conv_io_weight_win_33_232),
    .io_weight_win_33_233(conv_io_weight_win_33_233),
    .io_weight_win_33_234(conv_io_weight_win_33_234),
    .io_weight_win_33_235(conv_io_weight_win_33_235),
    .io_weight_win_33_236(conv_io_weight_win_33_236),
    .io_weight_win_33_237(conv_io_weight_win_33_237),
    .io_weight_win_33_238(conv_io_weight_win_33_238),
    .io_weight_win_33_239(conv_io_weight_win_33_239),
    .io_weight_win_33_240(conv_io_weight_win_33_240),
    .io_weight_win_33_241(conv_io_weight_win_33_241),
    .io_weight_win_33_242(conv_io_weight_win_33_242),
    .io_weight_win_33_243(conv_io_weight_win_33_243),
    .io_weight_win_33_244(conv_io_weight_win_33_244),
    .io_weight_win_33_245(conv_io_weight_win_33_245),
    .io_weight_win_33_246(conv_io_weight_win_33_246),
    .io_weight_win_33_247(conv_io_weight_win_33_247),
    .io_weight_win_33_248(conv_io_weight_win_33_248),
    .io_weight_win_33_249(conv_io_weight_win_33_249),
    .io_weight_win_33_250(conv_io_weight_win_33_250),
    .io_weight_win_33_251(conv_io_weight_win_33_251),
    .io_weight_win_33_252(conv_io_weight_win_33_252),
    .io_weight_win_33_253(conv_io_weight_win_33_253),
    .io_weight_win_33_254(conv_io_weight_win_33_254),
    .io_weight_win_33_255(conv_io_weight_win_33_255),
    .io_weight_win_33_256(conv_io_weight_win_33_256),
    .io_weight_win_33_257(conv_io_weight_win_33_257),
    .io_weight_win_33_258(conv_io_weight_win_33_258),
    .io_weight_win_33_259(conv_io_weight_win_33_259),
    .io_weight_win_33_260(conv_io_weight_win_33_260),
    .io_weight_win_33_261(conv_io_weight_win_33_261),
    .io_weight_win_33_262(conv_io_weight_win_33_262),
    .io_weight_win_33_263(conv_io_weight_win_33_263),
    .io_weight_win_33_264(conv_io_weight_win_33_264),
    .io_weight_win_33_265(conv_io_weight_win_33_265),
    .io_weight_win_33_266(conv_io_weight_win_33_266),
    .io_weight_win_33_267(conv_io_weight_win_33_267),
    .io_weight_win_33_268(conv_io_weight_win_33_268),
    .io_weight_win_33_269(conv_io_weight_win_33_269),
    .io_weight_win_33_270(conv_io_weight_win_33_270),
    .io_weight_win_33_271(conv_io_weight_win_33_271),
    .io_weight_win_33_272(conv_io_weight_win_33_272),
    .io_weight_win_33_273(conv_io_weight_win_33_273),
    .io_weight_win_33_274(conv_io_weight_win_33_274),
    .io_weight_win_33_275(conv_io_weight_win_33_275),
    .io_weight_win_33_276(conv_io_weight_win_33_276),
    .io_weight_win_33_277(conv_io_weight_win_33_277),
    .io_weight_win_33_278(conv_io_weight_win_33_278),
    .io_weight_win_33_279(conv_io_weight_win_33_279),
    .io_weight_win_33_280(conv_io_weight_win_33_280),
    .io_weight_win_33_281(conv_io_weight_win_33_281),
    .io_weight_win_33_282(conv_io_weight_win_33_282),
    .io_weight_win_33_283(conv_io_weight_win_33_283),
    .io_weight_win_33_284(conv_io_weight_win_33_284),
    .io_weight_win_33_285(conv_io_weight_win_33_285),
    .io_weight_win_33_286(conv_io_weight_win_33_286),
    .io_weight_win_33_287(conv_io_weight_win_33_287),
    .io_weight_win_33_288(conv_io_weight_win_33_288),
    .io_weight_win_33_289(conv_io_weight_win_33_289),
    .io_weight_win_33_290(conv_io_weight_win_33_290),
    .io_weight_win_33_291(conv_io_weight_win_33_291),
    .io_weight_win_33_292(conv_io_weight_win_33_292),
    .io_weight_win_33_293(conv_io_weight_win_33_293),
    .io_weight_win_33_294(conv_io_weight_win_33_294),
    .io_weight_win_33_295(conv_io_weight_win_33_295),
    .io_weight_win_33_296(conv_io_weight_win_33_296),
    .io_weight_win_33_297(conv_io_weight_win_33_297),
    .io_weight_win_33_298(conv_io_weight_win_33_298),
    .io_weight_win_33_299(conv_io_weight_win_33_299),
    .io_weight_win_33_300(conv_io_weight_win_33_300),
    .io_weight_win_33_301(conv_io_weight_win_33_301),
    .io_weight_win_33_302(conv_io_weight_win_33_302),
    .io_weight_win_33_303(conv_io_weight_win_33_303),
    .io_weight_win_33_304(conv_io_weight_win_33_304),
    .io_weight_win_33_305(conv_io_weight_win_33_305),
    .io_weight_win_33_306(conv_io_weight_win_33_306),
    .io_weight_win_33_307(conv_io_weight_win_33_307),
    .io_weight_win_33_308(conv_io_weight_win_33_308),
    .io_weight_win_33_309(conv_io_weight_win_33_309),
    .io_weight_win_33_310(conv_io_weight_win_33_310),
    .io_weight_win_33_311(conv_io_weight_win_33_311),
    .io_weight_win_33_312(conv_io_weight_win_33_312),
    .io_weight_win_33_313(conv_io_weight_win_33_313),
    .io_weight_win_33_314(conv_io_weight_win_33_314),
    .io_weight_win_33_315(conv_io_weight_win_33_315),
    .io_weight_win_33_316(conv_io_weight_win_33_316),
    .io_weight_win_33_317(conv_io_weight_win_33_317),
    .io_weight_win_33_318(conv_io_weight_win_33_318),
    .io_weight_win_33_319(conv_io_weight_win_33_319),
    .io_weight_win_33_320(conv_io_weight_win_33_320),
    .io_weight_win_33_321(conv_io_weight_win_33_321),
    .io_weight_win_33_322(conv_io_weight_win_33_322),
    .io_weight_win_33_323(conv_io_weight_win_33_323),
    .io_weight_win_33_324(conv_io_weight_win_33_324),
    .io_weight_win_33_325(conv_io_weight_win_33_325),
    .io_weight_win_33_326(conv_io_weight_win_33_326),
    .io_weight_win_33_327(conv_io_weight_win_33_327),
    .io_weight_win_33_328(conv_io_weight_win_33_328),
    .io_weight_win_33_329(conv_io_weight_win_33_329),
    .io_weight_win_33_330(conv_io_weight_win_33_330),
    .io_weight_win_33_331(conv_io_weight_win_33_331),
    .io_weight_win_33_332(conv_io_weight_win_33_332),
    .io_weight_win_33_333(conv_io_weight_win_33_333),
    .io_weight_win_33_334(conv_io_weight_win_33_334),
    .io_weight_win_33_335(conv_io_weight_win_33_335),
    .io_weight_win_33_336(conv_io_weight_win_33_336),
    .io_weight_win_33_337(conv_io_weight_win_33_337),
    .io_weight_win_33_338(conv_io_weight_win_33_338),
    .io_weight_win_33_339(conv_io_weight_win_33_339),
    .io_weight_win_33_340(conv_io_weight_win_33_340),
    .io_weight_win_33_341(conv_io_weight_win_33_341),
    .io_weight_win_33_342(conv_io_weight_win_33_342),
    .io_weight_win_33_343(conv_io_weight_win_33_343),
    .io_weight_win_33_344(conv_io_weight_win_33_344),
    .io_weight_win_33_345(conv_io_weight_win_33_345),
    .io_weight_win_33_346(conv_io_weight_win_33_346),
    .io_weight_win_33_347(conv_io_weight_win_33_347),
    .io_weight_win_33_348(conv_io_weight_win_33_348),
    .io_weight_win_33_349(conv_io_weight_win_33_349),
    .io_weight_win_33_350(conv_io_weight_win_33_350),
    .io_weight_win_33_351(conv_io_weight_win_33_351),
    .io_weight_win_33_352(conv_io_weight_win_33_352),
    .io_weight_win_33_353(conv_io_weight_win_33_353),
    .io_weight_win_33_354(conv_io_weight_win_33_354),
    .io_weight_win_33_355(conv_io_weight_win_33_355),
    .io_weight_win_33_356(conv_io_weight_win_33_356),
    .io_weight_win_33_357(conv_io_weight_win_33_357),
    .io_weight_win_33_358(conv_io_weight_win_33_358),
    .io_weight_win_33_359(conv_io_weight_win_33_359),
    .io_weight_win_33_360(conv_io_weight_win_33_360),
    .io_weight_win_33_361(conv_io_weight_win_33_361),
    .io_weight_win_33_362(conv_io_weight_win_33_362),
    .io_weight_win_33_363(conv_io_weight_win_33_363),
    .io_weight_win_33_364(conv_io_weight_win_33_364),
    .io_weight_win_33_365(conv_io_weight_win_33_365),
    .io_weight_win_33_366(conv_io_weight_win_33_366),
    .io_weight_win_33_367(conv_io_weight_win_33_367),
    .io_weight_win_33_368(conv_io_weight_win_33_368),
    .io_weight_win_33_369(conv_io_weight_win_33_369),
    .io_weight_win_33_370(conv_io_weight_win_33_370),
    .io_weight_win_33_371(conv_io_weight_win_33_371),
    .io_weight_win_33_372(conv_io_weight_win_33_372),
    .io_weight_win_33_373(conv_io_weight_win_33_373),
    .io_weight_win_33_374(conv_io_weight_win_33_374),
    .io_weight_win_33_375(conv_io_weight_win_33_375),
    .io_weight_win_33_376(conv_io_weight_win_33_376),
    .io_weight_win_33_377(conv_io_weight_win_33_377),
    .io_weight_win_33_378(conv_io_weight_win_33_378),
    .io_weight_win_33_379(conv_io_weight_win_33_379),
    .io_weight_win_33_380(conv_io_weight_win_33_380),
    .io_weight_win_33_381(conv_io_weight_win_33_381),
    .io_weight_win_33_382(conv_io_weight_win_33_382),
    .io_weight_win_33_383(conv_io_weight_win_33_383),
    .io_weight_win_33_384(conv_io_weight_win_33_384),
    .io_weight_win_33_385(conv_io_weight_win_33_385),
    .io_weight_win_33_386(conv_io_weight_win_33_386),
    .io_weight_win_33_387(conv_io_weight_win_33_387),
    .io_weight_win_33_388(conv_io_weight_win_33_388),
    .io_weight_win_33_389(conv_io_weight_win_33_389),
    .io_weight_win_33_390(conv_io_weight_win_33_390),
    .io_weight_win_33_391(conv_io_weight_win_33_391),
    .io_weight_win_33_392(conv_io_weight_win_33_392),
    .io_weight_win_33_393(conv_io_weight_win_33_393),
    .io_weight_win_33_394(conv_io_weight_win_33_394),
    .io_weight_win_33_395(conv_io_weight_win_33_395),
    .io_weight_win_33_396(conv_io_weight_win_33_396),
    .io_weight_win_33_397(conv_io_weight_win_33_397),
    .io_weight_win_33_398(conv_io_weight_win_33_398),
    .io_weight_win_33_399(conv_io_weight_win_33_399),
    .io_weight_win_33_400(conv_io_weight_win_33_400),
    .io_weight_win_33_401(conv_io_weight_win_33_401),
    .io_weight_win_33_402(conv_io_weight_win_33_402),
    .io_weight_win_33_403(conv_io_weight_win_33_403),
    .io_weight_win_33_404(conv_io_weight_win_33_404),
    .io_weight_win_33_405(conv_io_weight_win_33_405),
    .io_weight_win_33_406(conv_io_weight_win_33_406),
    .io_weight_win_33_407(conv_io_weight_win_33_407),
    .io_weight_win_33_408(conv_io_weight_win_33_408),
    .io_weight_win_33_409(conv_io_weight_win_33_409),
    .io_weight_win_33_410(conv_io_weight_win_33_410),
    .io_weight_win_33_411(conv_io_weight_win_33_411),
    .io_weight_win_33_412(conv_io_weight_win_33_412),
    .io_weight_win_33_413(conv_io_weight_win_33_413),
    .io_weight_win_33_414(conv_io_weight_win_33_414),
    .io_weight_win_33_415(conv_io_weight_win_33_415),
    .io_weight_win_33_416(conv_io_weight_win_33_416),
    .io_weight_win_33_417(conv_io_weight_win_33_417),
    .io_weight_win_33_418(conv_io_weight_win_33_418),
    .io_weight_win_33_419(conv_io_weight_win_33_419),
    .io_weight_win_33_420(conv_io_weight_win_33_420),
    .io_weight_win_33_421(conv_io_weight_win_33_421),
    .io_weight_win_33_422(conv_io_weight_win_33_422),
    .io_weight_win_33_423(conv_io_weight_win_33_423),
    .io_weight_win_33_424(conv_io_weight_win_33_424),
    .io_weight_win_33_425(conv_io_weight_win_33_425),
    .io_weight_win_33_426(conv_io_weight_win_33_426),
    .io_weight_win_33_427(conv_io_weight_win_33_427),
    .io_weight_win_33_428(conv_io_weight_win_33_428),
    .io_weight_win_33_429(conv_io_weight_win_33_429),
    .io_weight_win_33_430(conv_io_weight_win_33_430),
    .io_weight_win_33_431(conv_io_weight_win_33_431),
    .io_weight_win_33_432(conv_io_weight_win_33_432),
    .io_weight_win_33_433(conv_io_weight_win_33_433),
    .io_weight_win_33_434(conv_io_weight_win_33_434),
    .io_weight_win_33_435(conv_io_weight_win_33_435),
    .io_weight_win_33_436(conv_io_weight_win_33_436),
    .io_weight_win_33_437(conv_io_weight_win_33_437),
    .io_weight_win_33_438(conv_io_weight_win_33_438),
    .io_weight_win_33_439(conv_io_weight_win_33_439),
    .io_weight_win_33_440(conv_io_weight_win_33_440),
    .io_weight_win_33_441(conv_io_weight_win_33_441),
    .io_weight_win_33_442(conv_io_weight_win_33_442),
    .io_weight_win_33_443(conv_io_weight_win_33_443),
    .io_weight_win_33_444(conv_io_weight_win_33_444),
    .io_weight_win_33_445(conv_io_weight_win_33_445),
    .io_weight_win_33_446(conv_io_weight_win_33_446),
    .io_weight_win_33_447(conv_io_weight_win_33_447),
    .io_weight_win_33_448(conv_io_weight_win_33_448),
    .io_weight_win_33_449(conv_io_weight_win_33_449),
    .io_weight_win_33_450(conv_io_weight_win_33_450),
    .io_weight_win_33_451(conv_io_weight_win_33_451),
    .io_weight_win_33_452(conv_io_weight_win_33_452),
    .io_weight_win_33_453(conv_io_weight_win_33_453),
    .io_weight_win_33_454(conv_io_weight_win_33_454),
    .io_weight_win_33_455(conv_io_weight_win_33_455),
    .io_weight_win_33_456(conv_io_weight_win_33_456),
    .io_weight_win_33_457(conv_io_weight_win_33_457),
    .io_weight_win_33_458(conv_io_weight_win_33_458),
    .io_weight_win_33_459(conv_io_weight_win_33_459),
    .io_weight_win_33_460(conv_io_weight_win_33_460),
    .io_weight_win_33_461(conv_io_weight_win_33_461),
    .io_weight_win_33_462(conv_io_weight_win_33_462),
    .io_weight_win_33_463(conv_io_weight_win_33_463),
    .io_weight_win_33_464(conv_io_weight_win_33_464),
    .io_weight_win_33_465(conv_io_weight_win_33_465),
    .io_weight_win_33_466(conv_io_weight_win_33_466),
    .io_weight_win_33_467(conv_io_weight_win_33_467),
    .io_weight_win_33_468(conv_io_weight_win_33_468),
    .io_weight_win_33_469(conv_io_weight_win_33_469),
    .io_weight_win_33_470(conv_io_weight_win_33_470),
    .io_weight_win_33_471(conv_io_weight_win_33_471),
    .io_weight_win_33_472(conv_io_weight_win_33_472),
    .io_weight_win_33_473(conv_io_weight_win_33_473),
    .io_weight_win_33_474(conv_io_weight_win_33_474),
    .io_weight_win_33_475(conv_io_weight_win_33_475),
    .io_weight_win_33_476(conv_io_weight_win_33_476),
    .io_weight_win_33_477(conv_io_weight_win_33_477),
    .io_weight_win_33_478(conv_io_weight_win_33_478),
    .io_weight_win_33_479(conv_io_weight_win_33_479),
    .io_weight_win_33_480(conv_io_weight_win_33_480),
    .io_weight_win_33_481(conv_io_weight_win_33_481),
    .io_weight_win_33_482(conv_io_weight_win_33_482),
    .io_weight_win_33_483(conv_io_weight_win_33_483),
    .io_weight_win_33_484(conv_io_weight_win_33_484),
    .io_weight_win_33_485(conv_io_weight_win_33_485),
    .io_weight_win_33_486(conv_io_weight_win_33_486),
    .io_weight_win_33_487(conv_io_weight_win_33_487),
    .io_weight_win_33_488(conv_io_weight_win_33_488),
    .io_weight_win_33_489(conv_io_weight_win_33_489),
    .io_weight_win_33_490(conv_io_weight_win_33_490),
    .io_weight_win_33_491(conv_io_weight_win_33_491),
    .io_weight_win_33_492(conv_io_weight_win_33_492),
    .io_weight_win_33_493(conv_io_weight_win_33_493),
    .io_weight_win_33_494(conv_io_weight_win_33_494),
    .io_weight_win_33_495(conv_io_weight_win_33_495),
    .io_weight_win_33_496(conv_io_weight_win_33_496),
    .io_weight_win_33_497(conv_io_weight_win_33_497),
    .io_weight_win_33_498(conv_io_weight_win_33_498),
    .io_weight_win_33_499(conv_io_weight_win_33_499),
    .io_weight_win_33_500(conv_io_weight_win_33_500),
    .io_weight_win_33_501(conv_io_weight_win_33_501),
    .io_weight_win_33_502(conv_io_weight_win_33_502),
    .io_weight_win_33_503(conv_io_weight_win_33_503),
    .io_weight_win_33_504(conv_io_weight_win_33_504),
    .io_weight_win_33_505(conv_io_weight_win_33_505),
    .io_weight_win_33_506(conv_io_weight_win_33_506),
    .io_weight_win_33_507(conv_io_weight_win_33_507),
    .io_weight_win_33_508(conv_io_weight_win_33_508),
    .io_weight_win_33_509(conv_io_weight_win_33_509),
    .io_weight_win_33_510(conv_io_weight_win_33_510),
    .io_weight_win_33_511(conv_io_weight_win_33_511),
    .io_weight_win_33_512(conv_io_weight_win_33_512),
    .io_weight_win_33_513(conv_io_weight_win_33_513),
    .io_weight_win_33_514(conv_io_weight_win_33_514),
    .io_weight_win_33_515(conv_io_weight_win_33_515),
    .io_weight_win_33_516(conv_io_weight_win_33_516),
    .io_weight_win_33_517(conv_io_weight_win_33_517),
    .io_weight_win_33_518(conv_io_weight_win_33_518),
    .io_weight_win_33_519(conv_io_weight_win_33_519),
    .io_weight_win_33_520(conv_io_weight_win_33_520),
    .io_weight_win_33_521(conv_io_weight_win_33_521),
    .io_weight_win_33_522(conv_io_weight_win_33_522),
    .io_weight_win_33_523(conv_io_weight_win_33_523),
    .io_weight_win_33_524(conv_io_weight_win_33_524),
    .io_weight_win_33_525(conv_io_weight_win_33_525),
    .io_weight_win_33_526(conv_io_weight_win_33_526),
    .io_weight_win_33_527(conv_io_weight_win_33_527),
    .io_weight_win_33_528(conv_io_weight_win_33_528),
    .io_weight_win_33_529(conv_io_weight_win_33_529),
    .io_weight_win_33_530(conv_io_weight_win_33_530),
    .io_weight_win_33_531(conv_io_weight_win_33_531),
    .io_weight_win_33_532(conv_io_weight_win_33_532),
    .io_weight_win_33_533(conv_io_weight_win_33_533),
    .io_weight_win_33_534(conv_io_weight_win_33_534),
    .io_weight_win_33_535(conv_io_weight_win_33_535),
    .io_weight_win_33_536(conv_io_weight_win_33_536),
    .io_weight_win_33_537(conv_io_weight_win_33_537),
    .io_weight_win_33_538(conv_io_weight_win_33_538),
    .io_weight_win_33_539(conv_io_weight_win_33_539),
    .io_weight_win_33_540(conv_io_weight_win_33_540),
    .io_weight_win_33_541(conv_io_weight_win_33_541),
    .io_weight_win_33_542(conv_io_weight_win_33_542),
    .io_weight_win_33_543(conv_io_weight_win_33_543),
    .io_weight_win_33_544(conv_io_weight_win_33_544),
    .io_weight_win_33_545(conv_io_weight_win_33_545),
    .io_weight_win_33_546(conv_io_weight_win_33_546),
    .io_weight_win_33_547(conv_io_weight_win_33_547),
    .io_weight_win_33_548(conv_io_weight_win_33_548),
    .io_weight_win_33_549(conv_io_weight_win_33_549),
    .io_weight_win_33_550(conv_io_weight_win_33_550),
    .io_weight_win_33_551(conv_io_weight_win_33_551),
    .io_weight_win_33_552(conv_io_weight_win_33_552),
    .io_weight_win_33_553(conv_io_weight_win_33_553),
    .io_weight_win_33_554(conv_io_weight_win_33_554),
    .io_weight_win_33_555(conv_io_weight_win_33_555),
    .io_weight_win_33_556(conv_io_weight_win_33_556),
    .io_weight_win_33_557(conv_io_weight_win_33_557),
    .io_weight_win_33_558(conv_io_weight_win_33_558),
    .io_weight_win_33_559(conv_io_weight_win_33_559),
    .io_weight_win_33_560(conv_io_weight_win_33_560),
    .io_weight_win_33_561(conv_io_weight_win_33_561),
    .io_weight_win_33_562(conv_io_weight_win_33_562),
    .io_weight_win_33_563(conv_io_weight_win_33_563),
    .io_weight_win_33_564(conv_io_weight_win_33_564),
    .io_weight_win_33_565(conv_io_weight_win_33_565),
    .io_weight_win_33_566(conv_io_weight_win_33_566),
    .io_weight_win_33_567(conv_io_weight_win_33_567),
    .io_weight_win_33_568(conv_io_weight_win_33_568),
    .io_weight_win_33_569(conv_io_weight_win_33_569),
    .io_weight_win_33_570(conv_io_weight_win_33_570),
    .io_weight_win_33_571(conv_io_weight_win_33_571),
    .io_weight_win_33_572(conv_io_weight_win_33_572),
    .io_weight_win_33_573(conv_io_weight_win_33_573),
    .io_weight_win_33_574(conv_io_weight_win_33_574),
    .io_weight_win_33_575(conv_io_weight_win_33_575),
    .io_bias_data_0(conv_io_bias_data_0),
    .io_bias_data_1(conv_io_bias_data_1),
    .io_bias_data_2(conv_io_bias_data_2),
    .io_bias_data_3(conv_io_bias_data_3),
    .io_bias_data_4(conv_io_bias_data_4),
    .io_bias_data_5(conv_io_bias_data_5),
    .io_bias_data_6(conv_io_bias_data_6),
    .io_bias_data_7(conv_io_bias_data_7),
    .io_bias_valid(conv_io_bias_valid),
    .io_conv_o_0(conv_io_conv_o_0),
    .io_conv_o_1(conv_io_conv_o_1),
    .io_conv_o_2(conv_io_conv_o_2),
    .io_conv_o_3(conv_io_conv_o_3),
    .io_conv_o_4(conv_io_conv_o_4),
    .io_conv_o_5(conv_io_conv_o_5),
    .io_conv_o_6(conv_io_conv_o_6),
    .io_conv_o_7(conv_io_conv_o_7)
  );
  acc acc ( // @[acccel_top.scala 182:21]
    .clock(acc_clock),
    .reset(acc_reset),
    .io_prev_data_zero(acc_io_prev_data_zero),
    .io_curr_data_zero(acc_io_curr_data_zero),
    .io_read_en(acc_io_read_en),
    .io_write_en(acc_io_write_en),
    .io_read_addr(acc_io_read_addr),
    .io_write_addr(acc_io_write_addr),
    .io_curr_data_0(acc_io_curr_data_0),
    .io_curr_data_1(acc_io_curr_data_1),
    .io_curr_data_2(acc_io_curr_data_2),
    .io_curr_data_3(acc_io_curr_data_3),
    .io_curr_data_4(acc_io_curr_data_4),
    .io_curr_data_5(acc_io_curr_data_5),
    .io_curr_data_6(acc_io_curr_data_6),
    .io_curr_data_7(acc_io_curr_data_7),
    .io_acc_result_0(acc_io_acc_result_0),
    .io_acc_result_1(acc_io_acc_result_1),
    .io_acc_result_2(acc_io_acc_result_2),
    .io_acc_result_3(acc_io_acc_result_3),
    .io_acc_result_4(acc_io_acc_result_4),
    .io_acc_result_5(acc_io_acc_result_5),
    .io_acc_result_6(acc_io_acc_result_6),
    .io_acc_result_7(acc_io_acc_result_7)
  );
  quant quant ( // @[acccel_top.scala 195:23]
    .clock(quant_clock),
    .io_acc_result_0(quant_io_acc_result_0),
    .io_acc_result_1(quant_io_acc_result_1),
    .io_acc_result_2(quant_io_acc_result_2),
    .io_acc_result_3(quant_io_acc_result_3),
    .io_acc_result_4(quant_io_acc_result_4),
    .io_acc_result_5(quant_io_acc_result_5),
    .io_acc_result_6(quant_io_acc_result_6),
    .io_acc_result_7(quant_io_acc_result_7),
    .io_scale(quant_io_scale),
    .io_shift(quant_io_shift),
    .io_zero_point(quant_io_zero_point),
    .io_quant_result_0(quant_io_quant_result_0),
    .io_quant_result_1(quant_io_quant_result_1),
    .io_quant_result_2(quant_io_quant_result_2),
    .io_quant_result_3(quant_io_quant_result_3),
    .io_quant_result_4(quant_io_quant_result_4),
    .io_quant_result_5(quant_io_quant_result_5),
    .io_quant_result_6(quant_io_quant_result_6),
    .io_quant_result_7(quant_io_quant_result_7)
  );
  yolov8_maxpool_data_rwcontrol pool_ctrl ( // @[acccel_top.scala 234:27]
    .clock(pool_ctrl_clock),
    .reset(pool_ctrl_reset),
    .io_pool_enable(pool_ctrl_io_pool_enable),
    .io_zero_point(pool_ctrl_io_zero_point),
    .io_pool_finish(pool_ctrl_io_pool_finish),
    .io_pool_input_0(pool_ctrl_io_pool_input_0),
    .io_pool_input_1(pool_ctrl_io_pool_input_1),
    .io_pool_input_2(pool_ctrl_io_pool_input_2),
    .io_pool_input_3(pool_ctrl_io_pool_input_3),
    .io_pool_input_4(pool_ctrl_io_pool_input_4),
    .io_pool_input_5(pool_ctrl_io_pool_input_5),
    .io_pool_input_6(pool_ctrl_io_pool_input_6),
    .io_pool_input_7(pool_ctrl_io_pool_input_7),
    .io_last_data_of_row(pool_ctrl_io_last_data_of_row),
    .io_pool_outdata_valid(pool_ctrl_io_pool_outdata_valid),
    .io_ofm_write_addr(pool_ctrl_io_ofm_write_addr),
    .io_ofm_en_write(pool_ctrl_io_ofm_en_write),
    .io_ofm_read_addr(pool_ctrl_io_ofm_read_addr),
    .io_ofm_read_bundle(pool_ctrl_io_ofm_read_bundle),
    .io_row(pool_ctrl_io_row),
    .io_col(pool_ctrl_io_col)
  );
  MaxPool pool ( // @[acccel_top.scala 249:22]
    .clock(pool_clock),
    .reset(pool_reset),
    .io_input_0(pool_io_input_0),
    .io_input_1(pool_io_input_1),
    .io_input_2(pool_io_input_2),
    .io_input_3(pool_io_input_3),
    .io_input_4(pool_io_input_4),
    .io_input_5(pool_io_input_5),
    .io_input_6(pool_io_input_6),
    .io_input_7(pool_io_input_7),
    .io_last_data_of_row(pool_io_last_data_of_row),
    .io_output_0(pool_io_output_0),
    .io_output_1(pool_io_output_1),
    .io_output_2(pool_io_output_2),
    .io_output_3(pool_io_output_3),
    .io_output_4(pool_io_output_4),
    .io_output_5(pool_io_output_5),
    .io_output_6(pool_io_output_6),
    .io_output_7(pool_io_output_7),
    .io_outdata_valid(pool_io_outdata_valid)
  );
  BottleNeck_add bn_add ( // @[acccel_top.scala 276:24]
    .clock(bn_add_clock),
    .reset(bn_add_reset),
    .io_ifm_read_addr(bn_add_io_ifm_read_addr),
    .io_ifm_addr_read_sel(bn_add_io_ifm_addr_read_sel),
    .io_ifm_read_data_0(bn_add_io_ifm_read_data_0),
    .io_ifm_read_data_1(bn_add_io_ifm_read_data_1),
    .io_ifm_read_data_2(bn_add_io_ifm_read_data_2),
    .io_ifm_read_data_3(bn_add_io_ifm_read_data_3),
    .io_ifm_read_data_4(bn_add_io_ifm_read_data_4),
    .io_ifm_read_data_5(bn_add_io_ifm_read_data_5),
    .io_ifm_read_data_6(bn_add_io_ifm_read_data_6),
    .io_ifm_read_data_7(bn_add_io_ifm_read_data_7),
    .io_ofm_write_addr(bn_add_io_ofm_write_addr),
    .io_ofm_en_write(bn_add_io_ofm_en_write),
    .io_ofm_read_addr(bn_add_io_ofm_read_addr),
    .io_ofm_write_data(bn_add_io_ofm_write_data),
    .io_ofm_read_data(bn_add_io_ofm_read_data),
    .io_col(bn_add_io_col),
    .io_row(bn_add_io_row),
    .io_bottleneck_add_enable(bn_add_io_bottleneck_add_enable),
    .io_bottleneck_add_finish(bn_add_io_bottleneck_add_finish),
    .io_bn_add_in0_0(bn_add_io_bn_add_in0_0),
    .io_bn_add_in0_1(bn_add_io_bn_add_in0_1),
    .io_bn_add_in0_2(bn_add_io_bn_add_in0_2),
    .io_bn_add_in0_3(bn_add_io_bn_add_in0_3),
    .io_bn_add_in0_4(bn_add_io_bn_add_in0_4),
    .io_bn_add_in0_5(bn_add_io_bn_add_in0_5),
    .io_bn_add_in0_6(bn_add_io_bn_add_in0_6),
    .io_bn_add_in0_7(bn_add_io_bn_add_in0_7),
    .io_bn_add_in1_0(bn_add_io_bn_add_in1_0),
    .io_bn_add_in1_1(bn_add_io_bn_add_in1_1),
    .io_bn_add_in1_2(bn_add_io_bn_add_in1_2),
    .io_bn_add_in1_3(bn_add_io_bn_add_in1_3),
    .io_bn_add_in1_4(bn_add_io_bn_add_in1_4),
    .io_bn_add_in1_5(bn_add_io_bn_add_in1_5),
    .io_bn_add_in1_6(bn_add_io_bn_add_in1_6),
    .io_bn_add_in1_7(bn_add_io_bn_add_in1_7),
    .io_bn_add_result_0(bn_add_io_bn_add_result_0),
    .io_bn_add_result_1(bn_add_io_bn_add_result_1),
    .io_bn_add_result_2(bn_add_io_bn_add_result_2),
    .io_bn_add_result_3(bn_add_io_bn_add_result_3),
    .io_bn_add_result_4(bn_add_io_bn_add_result_4),
    .io_bn_add_result_5(bn_add_io_bn_add_result_5),
    .io_bn_add_result_6(bn_add_io_bn_add_result_6),
    .io_bn_add_result_7(bn_add_io_bn_add_result_7)
  );
  OfmBuffer ofm ( // @[acccel_top.scala 303:21]
    .clock(ofm_clock),
    .io_bram_write_addr(ofm_io_bram_write_addr),
    .io_bram_en_write(ofm_io_bram_en_write),
    .io_bram_read_addr(ofm_io_bram_read_addr),
    .io_ofm_store_bundle(ofm_io_ofm_store_bundle),
    .io_ofm_out_bundle(ofm_io_ofm_out_bundle)
  );
  assign io_ofm_out_bundle = ofm_io_ofm_out_bundle; // @[acccel_top.scala 222:31 308:20]
  assign io_pool_finish = pool_ctrl_io_pool_finish; // @[acccel_top.scala 231:25 237:17]
  assign io_bottleneck_add_finish = bn_add_io_bottleneck_add_finish; // @[acccel_top.scala 279:27 89:37]
  assign io_act_indata_0 = quant_io_quant_result_0; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_1 = quant_io_quant_result_1; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_2 = quant_io_quant_result_2; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_3 = quant_io_quant_result_3; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_4 = quant_io_quant_result_4; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_5 = quant_io_quant_result_5; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_6 = quant_io_quant_result_6; // @[acccel_top.scala 194:28 201:25]
  assign io_act_indata_7 = quant_io_quant_result_7; // @[acccel_top.scala 194:28 201:25]
  assign io_bn_add_in0_0 = bn_add_io_bn_add_in0_0; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_1 = bn_add_io_bn_add_in0_1; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_2 = bn_add_io_bn_add_in0_2; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_3 = bn_add_io_bn_add_in0_3; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_4 = bn_add_io_bn_add_in0_4; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_5 = bn_add_io_bn_add_in0_5; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_6 = bn_add_io_bn_add_in0_6; // @[acccel_top.scala 290:19]
  assign io_bn_add_in0_7 = bn_add_io_bn_add_in0_7; // @[acccel_top.scala 290:19]
  assign io_bn_add_in1_0 = bn_add_io_bn_add_in1_0; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_1 = bn_add_io_bn_add_in1_1; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_2 = bn_add_io_bn_add_in1_2; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_3 = bn_add_io_bn_add_in1_3; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_4 = bn_add_io_bn_add_in1_4; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_5 = bn_add_io_bn_add_in1_5; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_6 = bn_add_io_bn_add_in1_6; // @[acccel_top.scala 291:19]
  assign io_bn_add_in1_7 = bn_add_io_bn_add_in1_7; // @[acccel_top.scala 291:19]
  assign io_yolo_cls_data_before_compare = {conv_data_7,_ofm_conv_data_T_5}; // @[Cat.scala 33:92]
  assign ifm_buf_clock = clock;
  assign ifm_buf_reset = reset;
  assign ifm_buf_io_ifmbuf_bram_addr_read_s1 = _ifm_buf_io_ifmbuf_bram_addr_read_s1_T[10:0]; // @[acccel_top.scala 96:41]
  assign ifm_buf_io_ifmbuf_bram_addr_read_sel_s1 = bottleneck_work ? bn_add_ifm_addr_read_sel :
    io_ifmbuf_bram_addr_read_sel_s1; // @[acccel_top.scala 97:51]
  assign ifm_buf_io_ifmbuf_bram_addr_read_s2_singal = io_ifmbuf_bram_addr_read_s2_singal; // @[acccel_top.scala 98:48]
  assign ifm_buf_io_ifmbuf_bram_addr_read_s2_double = io_ifmbuf_bram_addr_read_s2_double; // @[acccel_top.scala 99:48]
  assign ifm_buf_io_bram_en_write = io_ifmbuf_bram_en_write; // @[acccel_top.scala 100:30]
  assign ifm_buf_io_upsample_enable = io_upsample_enable; // @[acccel_top.scala 103:32]
  assign ifm_buf_io_recv_done = io_recv_done; // @[acccel_top.scala 105:26]
  assign ifm_buf_io_buf_sel = io_ifmbuf_sel; // @[acccel_top.scala 101:24]
  assign ifm_buf_io_s_mod = io_s_mod; // @[acccel_top.scala 102:22]
  assign ifm_buf_io_col = io_col; // @[acccel_top.scala 104:20]
  assign ifm_buf_io_in_0 = io_ifm_in_0; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_1 = io_ifm_in_1; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_2 = io_ifm_in_2; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_3 = io_ifm_in_3; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_4 = io_ifm_in_4; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_5 = io_ifm_in_5; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_6 = io_ifm_in_6; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_in_7 = io_ifm_in_7; // @[acccel_top.scala 115:26]
  assign ifm_buf_io_pad_top = io_pad_top; // @[acccel_top.scala 106:24]
  assign ifm_buf_io_pad_bottom = io_pad_bottom; // @[acccel_top.scala 107:27]
  assign ifm_buf_io_pad_left_and_right = io_pad_left_and_right; // @[acccel_top.scala 108:35]
  assign ifm_buf_io_zero_pad_valid_s2 = io_zero_pad_valid_s2; // @[acccel_top.scala 109:34]
  assign ifm_buf_io_zero_pad_valid_s1 = io_zero_pad_valid_s1; // @[acccel_top.scala 110:34]
  assign ifm_buf_io_zero_point_in = io_zero_point_in; // @[acccel_top.scala 113:30]
  assign weight_buf_clock = clock;
  assign weight_buf_reset = reset;
  assign weight_buf_io_clear = io_weightbuf_waddr_clear; // @[acccel_top.scala 121:25]
  assign weight_buf_io_bram_write_en = io_weightbuf_bram_en_write; // @[acccel_top.scala 122:33]
  assign weight_buf_io_in_0 = io_weight_in_0; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_1 = io_weight_in_1; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_2 = io_weight_in_2; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_3 = io_weight_in_3; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_4 = io_weight_in_4; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_5 = io_weight_in_5; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_6 = io_weight_in_6; // @[acccel_top.scala 127:29]
  assign weight_buf_io_in_7 = io_weight_in_7; // @[acccel_top.scala 127:29]
  assign weight_buf_io_read_addr = io_weightbuf_read_addr; // @[acccel_top.scala 123:29]
  assign weight_buf_io_sel_when_kernal_is_1 = io_weight_sel; // @[acccel_top.scala 124:39]
  assign weight_buf_io_kernal = io_kernal; // @[acccel_top.scala 125:25]
  assign bias_buf_clock = clock;
  assign bias_buf_reset = reset;
  assign bias_buf_io_clear = io_biasbuf_waddr_clear; // @[acccel_top.scala 135:23]
  assign bias_buf_io_bias_in = io_bias_in; // @[acccel_top.scala 136:25]
  assign bias_buf_io_bram_addr_read = io_biasbuf_read_addr; // @[acccel_top.scala 137:32]
  assign bias_buf_io_bram_en_write = io_biasbuf_bram_en_write; // @[acccel_top.scala 138:31]
  assign sub_zero_clock = clock;
  assign sub_zero_reset = reset;
  assign sub_zero_io_zero_point = io_zero_point_in; // @[acccel_top.scala 145:28]
  assign sub_zero_io_data_in_0 = ifmstream_0[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_1 = ifmstream_0[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_2 = ifmstream_0[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_3 = ifmstream_0[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_4 = ifmstream_1[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_5 = ifmstream_1[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_6 = ifmstream_1[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_7 = ifmstream_1[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_8 = ifmstream_2[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_9 = ifmstream_2[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_10 = ifmstream_2[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_11 = ifmstream_2[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_12 = ifmstream_3[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_13 = ifmstream_3[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_14 = ifmstream_3[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_15 = ifmstream_3[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_16 = ifmstream_4[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_17 = ifmstream_4[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_18 = ifmstream_4[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_19 = ifmstream_4[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_20 = ifmstream_5[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_21 = ifmstream_5[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_22 = ifmstream_5[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_23 = ifmstream_5[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_24 = ifmstream_6[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_25 = ifmstream_6[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_26 = ifmstream_6[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_27 = ifmstream_6[31:24]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_28 = ifmstream_7[7:0]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_29 = ifmstream_7[15:8]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_30 = ifmstream_7[23:16]; // @[acccel_top.scala 148:59]
  assign sub_zero_io_data_in_31 = ifmstream_7[31:24]; // @[acccel_top.scala 148:59]
  assign line_buf_clock = clock;
  assign line_buf_reset = reset;
  assign line_buf_io_sel = io_sel; // @[acccel_top.scala 155:21]
  assign line_buf_io_s_mod = io_s_mod; // @[acccel_top.scala 157:23]
  assign line_buf_io_lineBuffer_i_data_0 = {ifmstream_sub_zp_0_hi,ifmstream_sub_zp_0_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_1 = {ifmstream_sub_zp_1_hi,ifmstream_sub_zp_1_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_2 = {ifmstream_sub_zp_2_hi,ifmstream_sub_zp_2_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_3 = {ifmstream_sub_zp_3_hi,ifmstream_sub_zp_3_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_4 = {ifmstream_sub_zp_4_hi,ifmstream_sub_zp_4_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_5 = {ifmstream_sub_zp_5_hi,ifmstream_sub_zp_5_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_6 = {ifmstream_sub_zp_6_hi,ifmstream_sub_zp_6_lo}; // @[Cat.scala 33:92]
  assign line_buf_io_lineBuffer_i_data_7 = {ifmstream_sub_zp_7_hi,ifmstream_sub_zp_7_lo}; // @[Cat.scala 33:92]
  assign conv_clock = clock;
  assign conv_io_ifm_win_33_0 = line_buf_io_lineBuffer_o_data_0; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_1 = line_buf_io_lineBuffer_o_data_1; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_2 = line_buf_io_lineBuffer_o_data_2; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_3 = line_buf_io_lineBuffer_o_data_3; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_4 = line_buf_io_lineBuffer_o_data_4; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_5 = line_buf_io_lineBuffer_o_data_5; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_6 = line_buf_io_lineBuffer_o_data_6; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_7 = line_buf_io_lineBuffer_o_data_7; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_8 = line_buf_io_lineBuffer_o_data_8; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_9 = line_buf_io_lineBuffer_o_data_9; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_10 = line_buf_io_lineBuffer_o_data_10; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_11 = line_buf_io_lineBuffer_o_data_11; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_12 = line_buf_io_lineBuffer_o_data_12; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_13 = line_buf_io_lineBuffer_o_data_13; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_14 = line_buf_io_lineBuffer_o_data_14; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_15 = line_buf_io_lineBuffer_o_data_15; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_16 = line_buf_io_lineBuffer_o_data_16; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_17 = line_buf_io_lineBuffer_o_data_17; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_18 = line_buf_io_lineBuffer_o_data_18; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_19 = line_buf_io_lineBuffer_o_data_19; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_20 = line_buf_io_lineBuffer_o_data_20; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_21 = line_buf_io_lineBuffer_o_data_21; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_22 = line_buf_io_lineBuffer_o_data_22; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_23 = line_buf_io_lineBuffer_o_data_23; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_24 = line_buf_io_lineBuffer_o_data_24; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_25 = line_buf_io_lineBuffer_o_data_25; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_26 = line_buf_io_lineBuffer_o_data_26; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_27 = line_buf_io_lineBuffer_o_data_27; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_28 = line_buf_io_lineBuffer_o_data_28; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_29 = line_buf_io_lineBuffer_o_data_29; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_30 = line_buf_io_lineBuffer_o_data_30; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_31 = line_buf_io_lineBuffer_o_data_31; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_32 = line_buf_io_lineBuffer_o_data_32; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_33 = line_buf_io_lineBuffer_o_data_33; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_34 = line_buf_io_lineBuffer_o_data_34; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_35 = line_buf_io_lineBuffer_o_data_35; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_36 = line_buf_io_lineBuffer_o_data_36; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_37 = line_buf_io_lineBuffer_o_data_37; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_38 = line_buf_io_lineBuffer_o_data_38; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_39 = line_buf_io_lineBuffer_o_data_39; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_40 = line_buf_io_lineBuffer_o_data_40; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_41 = line_buf_io_lineBuffer_o_data_41; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_42 = line_buf_io_lineBuffer_o_data_42; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_43 = line_buf_io_lineBuffer_o_data_43; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_44 = line_buf_io_lineBuffer_o_data_44; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_45 = line_buf_io_lineBuffer_o_data_45; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_46 = line_buf_io_lineBuffer_o_data_46; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_47 = line_buf_io_lineBuffer_o_data_47; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_48 = line_buf_io_lineBuffer_o_data_48; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_49 = line_buf_io_lineBuffer_o_data_49; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_50 = line_buf_io_lineBuffer_o_data_50; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_51 = line_buf_io_lineBuffer_o_data_51; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_52 = line_buf_io_lineBuffer_o_data_52; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_53 = line_buf_io_lineBuffer_o_data_53; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_54 = line_buf_io_lineBuffer_o_data_54; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_55 = line_buf_io_lineBuffer_o_data_55; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_56 = line_buf_io_lineBuffer_o_data_56; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_57 = line_buf_io_lineBuffer_o_data_57; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_58 = line_buf_io_lineBuffer_o_data_58; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_59 = line_buf_io_lineBuffer_o_data_59; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_60 = line_buf_io_lineBuffer_o_data_60; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_61 = line_buf_io_lineBuffer_o_data_61; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_62 = line_buf_io_lineBuffer_o_data_62; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_63 = line_buf_io_lineBuffer_o_data_63; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_64 = line_buf_io_lineBuffer_o_data_64; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_65 = line_buf_io_lineBuffer_o_data_65; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_66 = line_buf_io_lineBuffer_o_data_66; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_67 = line_buf_io_lineBuffer_o_data_67; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_68 = line_buf_io_lineBuffer_o_data_68; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_69 = line_buf_io_lineBuffer_o_data_69; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_70 = line_buf_io_lineBuffer_o_data_70; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_ifm_win_33_71 = line_buf_io_lineBuffer_o_data_71; // @[acccel_top.scala 153:23 162:20]
  assign conv_io_weight_win_33_0 = weight_win_0[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_1 = weight_win_0[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_2 = weight_win_0[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_3 = weight_win_0[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_4 = weight_win_0[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_5 = weight_win_0[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_6 = weight_win_0[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_7 = weight_win_0[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_8 = weight_win_0[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_9 = weight_win_1[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_10 = weight_win_1[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_11 = weight_win_1[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_12 = weight_win_1[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_13 = weight_win_1[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_14 = weight_win_1[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_15 = weight_win_1[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_16 = weight_win_1[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_17 = weight_win_1[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_18 = weight_win_2[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_19 = weight_win_2[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_20 = weight_win_2[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_21 = weight_win_2[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_22 = weight_win_2[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_23 = weight_win_2[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_24 = weight_win_2[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_25 = weight_win_2[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_26 = weight_win_2[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_27 = weight_win_3[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_28 = weight_win_3[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_29 = weight_win_3[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_30 = weight_win_3[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_31 = weight_win_3[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_32 = weight_win_3[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_33 = weight_win_3[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_34 = weight_win_3[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_35 = weight_win_3[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_36 = weight_win_4[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_37 = weight_win_4[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_38 = weight_win_4[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_39 = weight_win_4[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_40 = weight_win_4[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_41 = weight_win_4[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_42 = weight_win_4[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_43 = weight_win_4[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_44 = weight_win_4[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_45 = weight_win_5[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_46 = weight_win_5[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_47 = weight_win_5[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_48 = weight_win_5[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_49 = weight_win_5[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_50 = weight_win_5[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_51 = weight_win_5[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_52 = weight_win_5[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_53 = weight_win_5[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_54 = weight_win_6[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_55 = weight_win_6[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_56 = weight_win_6[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_57 = weight_win_6[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_58 = weight_win_6[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_59 = weight_win_6[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_60 = weight_win_6[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_61 = weight_win_6[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_62 = weight_win_6[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_63 = weight_win_7[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_64 = weight_win_7[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_65 = weight_win_7[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_66 = weight_win_7[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_67 = weight_win_7[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_68 = weight_win_7[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_69 = weight_win_7[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_70 = weight_win_7[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_71 = weight_win_7[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_72 = weight_win_8[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_73 = weight_win_8[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_74 = weight_win_8[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_75 = weight_win_8[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_76 = weight_win_8[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_77 = weight_win_8[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_78 = weight_win_8[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_79 = weight_win_8[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_80 = weight_win_8[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_81 = weight_win_9[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_82 = weight_win_9[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_83 = weight_win_9[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_84 = weight_win_9[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_85 = weight_win_9[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_86 = weight_win_9[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_87 = weight_win_9[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_88 = weight_win_9[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_89 = weight_win_9[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_90 = weight_win_10[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_91 = weight_win_10[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_92 = weight_win_10[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_93 = weight_win_10[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_94 = weight_win_10[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_95 = weight_win_10[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_96 = weight_win_10[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_97 = weight_win_10[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_98 = weight_win_10[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_99 = weight_win_11[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_100 = weight_win_11[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_101 = weight_win_11[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_102 = weight_win_11[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_103 = weight_win_11[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_104 = weight_win_11[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_105 = weight_win_11[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_106 = weight_win_11[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_107 = weight_win_11[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_108 = weight_win_12[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_109 = weight_win_12[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_110 = weight_win_12[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_111 = weight_win_12[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_112 = weight_win_12[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_113 = weight_win_12[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_114 = weight_win_12[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_115 = weight_win_12[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_116 = weight_win_12[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_117 = weight_win_13[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_118 = weight_win_13[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_119 = weight_win_13[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_120 = weight_win_13[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_121 = weight_win_13[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_122 = weight_win_13[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_123 = weight_win_13[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_124 = weight_win_13[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_125 = weight_win_13[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_126 = weight_win_14[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_127 = weight_win_14[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_128 = weight_win_14[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_129 = weight_win_14[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_130 = weight_win_14[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_131 = weight_win_14[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_132 = weight_win_14[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_133 = weight_win_14[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_134 = weight_win_14[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_135 = weight_win_15[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_136 = weight_win_15[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_137 = weight_win_15[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_138 = weight_win_15[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_139 = weight_win_15[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_140 = weight_win_15[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_141 = weight_win_15[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_142 = weight_win_15[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_143 = weight_win_15[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_144 = weight_win_16[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_145 = weight_win_16[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_146 = weight_win_16[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_147 = weight_win_16[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_148 = weight_win_16[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_149 = weight_win_16[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_150 = weight_win_16[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_151 = weight_win_16[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_152 = weight_win_16[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_153 = weight_win_17[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_154 = weight_win_17[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_155 = weight_win_17[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_156 = weight_win_17[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_157 = weight_win_17[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_158 = weight_win_17[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_159 = weight_win_17[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_160 = weight_win_17[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_161 = weight_win_17[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_162 = weight_win_18[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_163 = weight_win_18[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_164 = weight_win_18[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_165 = weight_win_18[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_166 = weight_win_18[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_167 = weight_win_18[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_168 = weight_win_18[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_169 = weight_win_18[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_170 = weight_win_18[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_171 = weight_win_19[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_172 = weight_win_19[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_173 = weight_win_19[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_174 = weight_win_19[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_175 = weight_win_19[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_176 = weight_win_19[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_177 = weight_win_19[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_178 = weight_win_19[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_179 = weight_win_19[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_180 = weight_win_20[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_181 = weight_win_20[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_182 = weight_win_20[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_183 = weight_win_20[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_184 = weight_win_20[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_185 = weight_win_20[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_186 = weight_win_20[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_187 = weight_win_20[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_188 = weight_win_20[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_189 = weight_win_21[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_190 = weight_win_21[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_191 = weight_win_21[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_192 = weight_win_21[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_193 = weight_win_21[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_194 = weight_win_21[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_195 = weight_win_21[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_196 = weight_win_21[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_197 = weight_win_21[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_198 = weight_win_22[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_199 = weight_win_22[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_200 = weight_win_22[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_201 = weight_win_22[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_202 = weight_win_22[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_203 = weight_win_22[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_204 = weight_win_22[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_205 = weight_win_22[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_206 = weight_win_22[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_207 = weight_win_23[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_208 = weight_win_23[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_209 = weight_win_23[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_210 = weight_win_23[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_211 = weight_win_23[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_212 = weight_win_23[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_213 = weight_win_23[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_214 = weight_win_23[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_215 = weight_win_23[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_216 = weight_win_24[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_217 = weight_win_24[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_218 = weight_win_24[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_219 = weight_win_24[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_220 = weight_win_24[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_221 = weight_win_24[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_222 = weight_win_24[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_223 = weight_win_24[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_224 = weight_win_24[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_225 = weight_win_25[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_226 = weight_win_25[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_227 = weight_win_25[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_228 = weight_win_25[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_229 = weight_win_25[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_230 = weight_win_25[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_231 = weight_win_25[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_232 = weight_win_25[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_233 = weight_win_25[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_234 = weight_win_26[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_235 = weight_win_26[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_236 = weight_win_26[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_237 = weight_win_26[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_238 = weight_win_26[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_239 = weight_win_26[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_240 = weight_win_26[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_241 = weight_win_26[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_242 = weight_win_26[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_243 = weight_win_27[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_244 = weight_win_27[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_245 = weight_win_27[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_246 = weight_win_27[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_247 = weight_win_27[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_248 = weight_win_27[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_249 = weight_win_27[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_250 = weight_win_27[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_251 = weight_win_27[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_252 = weight_win_28[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_253 = weight_win_28[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_254 = weight_win_28[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_255 = weight_win_28[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_256 = weight_win_28[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_257 = weight_win_28[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_258 = weight_win_28[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_259 = weight_win_28[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_260 = weight_win_28[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_261 = weight_win_29[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_262 = weight_win_29[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_263 = weight_win_29[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_264 = weight_win_29[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_265 = weight_win_29[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_266 = weight_win_29[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_267 = weight_win_29[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_268 = weight_win_29[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_269 = weight_win_29[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_270 = weight_win_30[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_271 = weight_win_30[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_272 = weight_win_30[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_273 = weight_win_30[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_274 = weight_win_30[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_275 = weight_win_30[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_276 = weight_win_30[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_277 = weight_win_30[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_278 = weight_win_30[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_279 = weight_win_31[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_280 = weight_win_31[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_281 = weight_win_31[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_282 = weight_win_31[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_283 = weight_win_31[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_284 = weight_win_31[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_285 = weight_win_31[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_286 = weight_win_31[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_287 = weight_win_31[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_288 = weight_win_32[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_289 = weight_win_32[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_290 = weight_win_32[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_291 = weight_win_32[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_292 = weight_win_32[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_293 = weight_win_32[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_294 = weight_win_32[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_295 = weight_win_32[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_296 = weight_win_32[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_297 = weight_win_33[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_298 = weight_win_33[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_299 = weight_win_33[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_300 = weight_win_33[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_301 = weight_win_33[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_302 = weight_win_33[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_303 = weight_win_33[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_304 = weight_win_33[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_305 = weight_win_33[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_306 = weight_win_34[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_307 = weight_win_34[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_308 = weight_win_34[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_309 = weight_win_34[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_310 = weight_win_34[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_311 = weight_win_34[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_312 = weight_win_34[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_313 = weight_win_34[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_314 = weight_win_34[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_315 = weight_win_35[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_316 = weight_win_35[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_317 = weight_win_35[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_318 = weight_win_35[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_319 = weight_win_35[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_320 = weight_win_35[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_321 = weight_win_35[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_322 = weight_win_35[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_323 = weight_win_35[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_324 = weight_win_36[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_325 = weight_win_36[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_326 = weight_win_36[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_327 = weight_win_36[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_328 = weight_win_36[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_329 = weight_win_36[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_330 = weight_win_36[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_331 = weight_win_36[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_332 = weight_win_36[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_333 = weight_win_37[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_334 = weight_win_37[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_335 = weight_win_37[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_336 = weight_win_37[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_337 = weight_win_37[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_338 = weight_win_37[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_339 = weight_win_37[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_340 = weight_win_37[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_341 = weight_win_37[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_342 = weight_win_38[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_343 = weight_win_38[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_344 = weight_win_38[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_345 = weight_win_38[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_346 = weight_win_38[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_347 = weight_win_38[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_348 = weight_win_38[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_349 = weight_win_38[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_350 = weight_win_38[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_351 = weight_win_39[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_352 = weight_win_39[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_353 = weight_win_39[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_354 = weight_win_39[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_355 = weight_win_39[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_356 = weight_win_39[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_357 = weight_win_39[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_358 = weight_win_39[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_359 = weight_win_39[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_360 = weight_win_40[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_361 = weight_win_40[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_362 = weight_win_40[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_363 = weight_win_40[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_364 = weight_win_40[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_365 = weight_win_40[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_366 = weight_win_40[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_367 = weight_win_40[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_368 = weight_win_40[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_369 = weight_win_41[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_370 = weight_win_41[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_371 = weight_win_41[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_372 = weight_win_41[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_373 = weight_win_41[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_374 = weight_win_41[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_375 = weight_win_41[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_376 = weight_win_41[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_377 = weight_win_41[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_378 = weight_win_42[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_379 = weight_win_42[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_380 = weight_win_42[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_381 = weight_win_42[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_382 = weight_win_42[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_383 = weight_win_42[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_384 = weight_win_42[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_385 = weight_win_42[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_386 = weight_win_42[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_387 = weight_win_43[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_388 = weight_win_43[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_389 = weight_win_43[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_390 = weight_win_43[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_391 = weight_win_43[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_392 = weight_win_43[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_393 = weight_win_43[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_394 = weight_win_43[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_395 = weight_win_43[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_396 = weight_win_44[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_397 = weight_win_44[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_398 = weight_win_44[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_399 = weight_win_44[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_400 = weight_win_44[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_401 = weight_win_44[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_402 = weight_win_44[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_403 = weight_win_44[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_404 = weight_win_44[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_405 = weight_win_45[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_406 = weight_win_45[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_407 = weight_win_45[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_408 = weight_win_45[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_409 = weight_win_45[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_410 = weight_win_45[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_411 = weight_win_45[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_412 = weight_win_45[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_413 = weight_win_45[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_414 = weight_win_46[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_415 = weight_win_46[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_416 = weight_win_46[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_417 = weight_win_46[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_418 = weight_win_46[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_419 = weight_win_46[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_420 = weight_win_46[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_421 = weight_win_46[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_422 = weight_win_46[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_423 = weight_win_47[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_424 = weight_win_47[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_425 = weight_win_47[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_426 = weight_win_47[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_427 = weight_win_47[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_428 = weight_win_47[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_429 = weight_win_47[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_430 = weight_win_47[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_431 = weight_win_47[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_432 = weight_win_48[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_433 = weight_win_48[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_434 = weight_win_48[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_435 = weight_win_48[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_436 = weight_win_48[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_437 = weight_win_48[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_438 = weight_win_48[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_439 = weight_win_48[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_440 = weight_win_48[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_441 = weight_win_49[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_442 = weight_win_49[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_443 = weight_win_49[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_444 = weight_win_49[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_445 = weight_win_49[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_446 = weight_win_49[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_447 = weight_win_49[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_448 = weight_win_49[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_449 = weight_win_49[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_450 = weight_win_50[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_451 = weight_win_50[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_452 = weight_win_50[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_453 = weight_win_50[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_454 = weight_win_50[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_455 = weight_win_50[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_456 = weight_win_50[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_457 = weight_win_50[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_458 = weight_win_50[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_459 = weight_win_51[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_460 = weight_win_51[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_461 = weight_win_51[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_462 = weight_win_51[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_463 = weight_win_51[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_464 = weight_win_51[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_465 = weight_win_51[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_466 = weight_win_51[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_467 = weight_win_51[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_468 = weight_win_52[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_469 = weight_win_52[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_470 = weight_win_52[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_471 = weight_win_52[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_472 = weight_win_52[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_473 = weight_win_52[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_474 = weight_win_52[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_475 = weight_win_52[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_476 = weight_win_52[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_477 = weight_win_53[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_478 = weight_win_53[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_479 = weight_win_53[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_480 = weight_win_53[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_481 = weight_win_53[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_482 = weight_win_53[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_483 = weight_win_53[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_484 = weight_win_53[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_485 = weight_win_53[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_486 = weight_win_54[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_487 = weight_win_54[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_488 = weight_win_54[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_489 = weight_win_54[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_490 = weight_win_54[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_491 = weight_win_54[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_492 = weight_win_54[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_493 = weight_win_54[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_494 = weight_win_54[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_495 = weight_win_55[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_496 = weight_win_55[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_497 = weight_win_55[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_498 = weight_win_55[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_499 = weight_win_55[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_500 = weight_win_55[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_501 = weight_win_55[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_502 = weight_win_55[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_503 = weight_win_55[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_504 = weight_win_56[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_505 = weight_win_56[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_506 = weight_win_56[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_507 = weight_win_56[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_508 = weight_win_56[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_509 = weight_win_56[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_510 = weight_win_56[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_511 = weight_win_56[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_512 = weight_win_56[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_513 = weight_win_57[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_514 = weight_win_57[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_515 = weight_win_57[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_516 = weight_win_57[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_517 = weight_win_57[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_518 = weight_win_57[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_519 = weight_win_57[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_520 = weight_win_57[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_521 = weight_win_57[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_522 = weight_win_58[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_523 = weight_win_58[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_524 = weight_win_58[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_525 = weight_win_58[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_526 = weight_win_58[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_527 = weight_win_58[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_528 = weight_win_58[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_529 = weight_win_58[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_530 = weight_win_58[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_531 = weight_win_59[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_532 = weight_win_59[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_533 = weight_win_59[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_534 = weight_win_59[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_535 = weight_win_59[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_536 = weight_win_59[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_537 = weight_win_59[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_538 = weight_win_59[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_539 = weight_win_59[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_540 = weight_win_60[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_541 = weight_win_60[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_542 = weight_win_60[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_543 = weight_win_60[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_544 = weight_win_60[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_545 = weight_win_60[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_546 = weight_win_60[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_547 = weight_win_60[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_548 = weight_win_60[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_549 = weight_win_61[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_550 = weight_win_61[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_551 = weight_win_61[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_552 = weight_win_61[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_553 = weight_win_61[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_554 = weight_win_61[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_555 = weight_win_61[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_556 = weight_win_61[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_557 = weight_win_61[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_558 = weight_win_62[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_559 = weight_win_62[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_560 = weight_win_62[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_561 = weight_win_62[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_562 = weight_win_62[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_563 = weight_win_62[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_564 = weight_win_62[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_565 = weight_win_62[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_566 = weight_win_62[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_567 = weight_win_63[7:0]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_568 = weight_win_63[15:8]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_569 = weight_win_63[23:16]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_570 = weight_win_63[31:24]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_571 = weight_win_63[39:32]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_572 = weight_win_63[47:40]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_573 = weight_win_63[55:48]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_574 = weight_win_63[63:56]; // @[acccel_top.scala 173:62]
  assign conv_io_weight_win_33_575 = weight_win_63[71:64]; // @[acccel_top.scala 173:62]
  assign conv_io_bias_data_0 = bias_buf_io_bias_data_0; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_1 = bias_buf_io_bias_data_1; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_2 = bias_buf_io_bias_data_2; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_3 = bias_buf_io_bias_data_3; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_4 = bias_buf_io_bias_data_4; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_5 = bias_buf_io_bias_data_5; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_6 = bias_buf_io_bias_data_6; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_data_7 = bias_buf_io_bias_data_7; // @[acccel_top.scala 133:20 140:17]
  assign conv_io_bias_valid = io_bias_valid; // @[acccel_top.scala 167:24]
  assign acc_clock = clock;
  assign acc_reset = reset;
  assign acc_io_prev_data_zero = io_acc_prev_data_zero; // @[acccel_top.scala 183:27]
  assign acc_io_curr_data_zero = io_acc_curr_data_zero; // @[acccel_top.scala 184:27]
  assign acc_io_read_en = io_acc_read_en; // @[acccel_top.scala 185:20]
  assign acc_io_write_en = io_acc_write_en; // @[acccel_top.scala 186:21]
  assign acc_io_read_addr = io_acc_read_addr; // @[acccel_top.scala 187:22]
  assign acc_io_write_addr = io_acc_write_addr; // @[acccel_top.scala 188:23]
  assign acc_io_curr_data_0 = conv_io_conv_o_0; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_1 = conv_io_conv_o_1; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_2 = conv_io_conv_o_2; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_3 = conv_io_conv_o_3; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_4 = conv_io_conv_o_4; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_5 = conv_io_conv_o_5; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_6 = conv_io_conv_o_6; // @[acccel_top.scala 165:29 178:26]
  assign acc_io_curr_data_7 = conv_io_conv_o_7; // @[acccel_top.scala 165:29 178:26]
  assign quant_clock = clock;
  assign quant_io_acc_result_0 = acc_io_acc_result_0; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_1 = acc_io_acc_result_1; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_2 = acc_io_acc_result_2; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_3 = acc_io_acc_result_3; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_4 = acc_io_acc_result_4; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_5 = acc_io_acc_result_5; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_6 = acc_io_acc_result_6; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_acc_result_7 = acc_io_acc_result_7; // @[acccel_top.scala 181:26 191:23]
  assign quant_io_scale = io_scale; // @[acccel_top.scala 196:20]
  assign quant_io_shift = io_shift; // @[acccel_top.scala 197:20]
  assign quant_io_zero_point = io_zero_point_out; // @[acccel_top.scala 198:25]
  assign pool_ctrl_clock = clock;
  assign pool_ctrl_reset = reset;
  assign pool_ctrl_io_pool_enable = io_pool_enable; // @[acccel_top.scala 235:30]
  assign pool_ctrl_io_zero_point = io_zero_point_A_act; // @[acccel_top.scala 236:29]
  assign pool_ctrl_io_pool_outdata_valid = pool_io_outdata_valid; // @[acccel_top.scala 251:37]
  assign pool_ctrl_io_ofm_read_bundle = ofm_io_ofm_out_bundle; // @[acccel_top.scala 222:31 308:20]
  assign pool_ctrl_io_row = io_row; // @[acccel_top.scala 243:22]
  assign pool_ctrl_io_col = io_col; // @[acccel_top.scala 244:22]
  assign pool_clock = clock;
  assign pool_reset = reset;
  assign pool_io_input_0 = pool_ctrl_io_pool_input_0; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_1 = pool_ctrl_io_pool_input_1; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_2 = pool_ctrl_io_pool_input_2; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_3 = pool_ctrl_io_pool_input_3; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_4 = pool_ctrl_io_pool_input_4; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_5 = pool_ctrl_io_pool_input_5; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_6 = pool_ctrl_io_pool_input_6; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_input_7 = pool_ctrl_io_pool_input_7; // @[acccel_top.scala 229:26 246:16]
  assign pool_io_last_data_of_row = pool_ctrl_io_last_data_of_row; // @[acccel_top.scala 250:30]
  assign bn_add_clock = clock;
  assign bn_add_reset = reset;
  assign bn_add_io_ifm_read_data_0 = ifmstream_0[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_1 = ifmstream_1[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_2 = ifmstream_2[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_3 = ifmstream_3[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_4 = ifmstream_4[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_5 = ifmstream_5[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_6 = ifmstream_6[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ifm_read_data_7 = ifmstream_7[7:0]; // @[acccel_top.scala 273:47]
  assign bn_add_io_ofm_read_data = ofm_io_ofm_out_bundle; // @[acccel_top.scala 222:31 308:20]
  assign bn_add_io_col = io_col; // @[acccel_top.scala 277:19]
  assign bn_add_io_row = io_row; // @[acccel_top.scala 278:19]
  assign bn_add_io_bottleneck_add_enable = io_bottleneck_add_enable; // @[acccel_top.scala 280:37]
  assign bn_add_io_bn_add_result_0 = io_bn_add_result_0; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_1 = io_bn_add_result_1; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_2 = io_bn_add_result_2; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_3 = io_bn_add_result_3; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_4 = io_bn_add_result_4; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_5 = io_bn_add_result_5; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_6 = io_bn_add_result_6; // @[acccel_top.scala 292:29]
  assign bn_add_io_bn_add_result_7 = io_bn_add_result_7; // @[acccel_top.scala 292:29]
  assign ofm_clock = clock;
  assign ofm_io_bram_write_addr = pool_work ? pool_ofm_write_addr : _ofm_write_addr_T; // @[acccel_top.scala 298:29]
  assign ofm_io_bram_en_write = pool_work ? pool_ofm_en_write : _ofm_en_write_T; // @[acccel_top.scala 299:27]
  assign ofm_io_bram_read_addr = ofm_read_addr[11:0]; // @[acccel_top.scala 305:27]
  assign ofm_io_ofm_store_bundle = pool_work ? pool_data_bundle : _ofm_store_bundle_T; // @[acccel_top.scala 301:31]
  always @(posedge clock) begin
    if (reset) begin // @[acccel_top.scala 88:34]
      bottleneck_work <= 1'h0; // @[acccel_top.scala 88:34]
    end else begin
      bottleneck_work <= _bottleneck_work_T_1 | _bottleneck_work_T_4; // @[acccel_top.scala 90:21]
    end
    if (reset) begin // @[utils.scala 10:17]
      bottleneck_work_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      bottleneck_work_REG <= io_bottleneck_add_enable; // @[utils.scala 10:17]
    end
    if (reset) begin // @[utils.scala 10:17]
      bottleneck_work_REG_1 <= 1'h0; // @[utils.scala 10:17]
    end else begin
      bottleneck_work_REG_1 <= bottleneck_add_finish; // @[utils.scala 10:17]
    end
    if (reset) begin // @[acccel_top.scala 294:28]
      pool_work <= 1'h0; // @[acccel_top.scala 294:28]
    end else begin
      pool_work <= _pool_work_T_1 | _pool_work_T_4; // @[acccel_top.scala 295:15]
    end
    if (reset) begin // @[utils.scala 10:17]
      pool_work_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      pool_work_REG <= io_pool_enable; // @[utils.scala 10:17]
    end
    if (reset) begin // @[utils.scala 10:17]
      pool_work_REG_1 <= 1'h0; // @[utils.scala 10:17]
    end else begin
      pool_work_REG_1 <= pool_finish; // @[utils.scala 10:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bottleneck_work = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  bottleneck_work_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  bottleneck_work_REG_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pool_work = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  pool_work_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  pool_work_REG_1 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module compare_8_cell(
  input         clock,
  input         reset,
  input         io_yolo_layer_finish,
  input  [63:0] io_data,
  output [7:0]  io_max_data,
  output [2:0]  io_max_index
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] data_0 = io_data[7:0]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_1 = io_data[15:8]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_2 = io_data[23:16]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_3 = io_data[31:24]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_4 = io_data[39:32]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_5 = io_data[47:40]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_6 = io_data[55:48]; // @[yolo_layer.scala 399:31]
  wire [7:0] data_7 = io_data[63:56]; // @[yolo_layer.scala 399:31]
  wire  _T_1 = reset | io_yolo_layer_finish; // @[yolo_layer.scala 401:32]
  reg [7:0] temp0_data_0; // @[yolo_layer.scala 403:49]
  reg [7:0] temp0_data_1; // @[yolo_layer.scala 403:49]
  reg [7:0] temp0_data_2; // @[yolo_layer.scala 403:49]
  reg [7:0] temp0_data_3; // @[yolo_layer.scala 403:49]
  reg [2:0] temp0_index_0; // @[yolo_layer.scala 404:50]
  reg [2:0] temp0_index_1; // @[yolo_layer.scala 404:50]
  reg [2:0] temp0_index_2; // @[yolo_layer.scala 404:50]
  reg [2:0] temp0_index_3; // @[yolo_layer.scala 404:50]
  wire  select0_0 = data_0 > data_1; // @[yolo_layer.scala 409:47]
  wire  _temp0_index_0_T = select0_0 ? 1'h0 : 1'h1; // @[yolo_layer.scala 412:38]
  wire  select0_1 = data_2 > data_3; // @[yolo_layer.scala 409:47]
  wire [1:0] _temp0_index_1_T = select0_1 ? 2'h2 : 2'h3; // @[yolo_layer.scala 412:38]
  wire  select0_2 = data_4 > data_5; // @[yolo_layer.scala 409:47]
  wire  select0_3 = data_6 > data_7; // @[yolo_layer.scala 409:47]
  reg [7:0] temp1_data_0; // @[yolo_layer.scala 416:49]
  reg [7:0] temp1_data_1; // @[yolo_layer.scala 416:49]
  reg [2:0] temp1_index_0; // @[yolo_layer.scala 417:50]
  reg [2:0] temp1_index_1; // @[yolo_layer.scala 417:50]
  wire  select1_0 = temp0_data_0 > temp0_data_1; // @[yolo_layer.scala 422:53]
  wire  select1_1 = temp0_data_2 > temp0_data_3; // @[yolo_layer.scala 422:53]
  reg [7:0] temp2_data_0; // @[yolo_layer.scala 429:49]
  reg [2:0] temp2_index_0; // @[yolo_layer.scala 430:50]
  wire  select2_0 = temp1_data_0 > temp1_data_1; // @[yolo_layer.scala 435:53]
  assign io_max_data = temp2_data_0; // @[yolo_layer.scala 440:25]
  assign io_max_index = temp2_index_0; // @[yolo_layer.scala 441:26]
  always @(posedge clock) begin
    if (_T_1) begin // @[yolo_layer.scala 403:49]
      temp0_data_0 <= 8'h0; // @[yolo_layer.scala 403:49]
    end else if (select0_0) begin // @[yolo_layer.scala 411:37]
      temp0_data_0 <= data_0;
    end else begin
      temp0_data_0 <= data_1;
    end
    if (_T_1) begin // @[yolo_layer.scala 403:49]
      temp0_data_1 <= 8'h0; // @[yolo_layer.scala 403:49]
    end else if (select0_1) begin // @[yolo_layer.scala 411:37]
      temp0_data_1 <= data_2;
    end else begin
      temp0_data_1 <= data_3;
    end
    if (_T_1) begin // @[yolo_layer.scala 403:49]
      temp0_data_2 <= 8'h0; // @[yolo_layer.scala 403:49]
    end else if (select0_2) begin // @[yolo_layer.scala 411:37]
      temp0_data_2 <= data_4;
    end else begin
      temp0_data_2 <= data_5;
    end
    if (_T_1) begin // @[yolo_layer.scala 403:49]
      temp0_data_3 <= 8'h0; // @[yolo_layer.scala 403:49]
    end else if (select0_3) begin // @[yolo_layer.scala 411:37]
      temp0_data_3 <= data_6;
    end else begin
      temp0_data_3 <= data_7;
    end
    if (_T_1) begin // @[yolo_layer.scala 404:50]
      temp0_index_0 <= 3'h0; // @[yolo_layer.scala 404:50]
    end else begin
      temp0_index_0 <= {{2'd0}, _temp0_index_0_T}; // @[yolo_layer.scala 412:32]
    end
    if (_T_1) begin // @[yolo_layer.scala 404:50]
      temp0_index_1 <= 3'h0; // @[yolo_layer.scala 404:50]
    end else begin
      temp0_index_1 <= {{1'd0}, _temp0_index_1_T}; // @[yolo_layer.scala 412:32]
    end
    if (_T_1) begin // @[yolo_layer.scala 404:50]
      temp0_index_2 <= 3'h0; // @[yolo_layer.scala 404:50]
    end else if (select0_2) begin // @[yolo_layer.scala 412:38]
      temp0_index_2 <= 3'h4;
    end else begin
      temp0_index_2 <= 3'h5;
    end
    if (_T_1) begin // @[yolo_layer.scala 404:50]
      temp0_index_3 <= 3'h0; // @[yolo_layer.scala 404:50]
    end else if (select0_3) begin // @[yolo_layer.scala 412:38]
      temp0_index_3 <= 3'h6;
    end else begin
      temp0_index_3 <= 3'h7;
    end
    if (_T_1) begin // @[yolo_layer.scala 416:49]
      temp1_data_0 <= 8'h0; // @[yolo_layer.scala 416:49]
    end else if (select1_0) begin // @[yolo_layer.scala 424:37]
      temp1_data_0 <= temp0_data_0;
    end else begin
      temp1_data_0 <= temp0_data_1;
    end
    if (_T_1) begin // @[yolo_layer.scala 416:49]
      temp1_data_1 <= 8'h0; // @[yolo_layer.scala 416:49]
    end else if (select1_1) begin // @[yolo_layer.scala 424:37]
      temp1_data_1 <= temp0_data_2;
    end else begin
      temp1_data_1 <= temp0_data_3;
    end
    if (_T_1) begin // @[yolo_layer.scala 417:50]
      temp1_index_0 <= 3'h0; // @[yolo_layer.scala 417:50]
    end else if (select1_0) begin // @[yolo_layer.scala 425:38]
      temp1_index_0 <= temp0_index_0;
    end else begin
      temp1_index_0 <= temp0_index_1;
    end
    if (_T_1) begin // @[yolo_layer.scala 417:50]
      temp1_index_1 <= 3'h0; // @[yolo_layer.scala 417:50]
    end else if (select1_1) begin // @[yolo_layer.scala 425:38]
      temp1_index_1 <= temp0_index_2;
    end else begin
      temp1_index_1 <= temp0_index_3;
    end
    if (_T_1) begin // @[yolo_layer.scala 429:49]
      temp2_data_0 <= 8'h0; // @[yolo_layer.scala 429:49]
    end else if (select2_0) begin // @[yolo_layer.scala 437:37]
      temp2_data_0 <= temp1_data_0;
    end else begin
      temp2_data_0 <= temp1_data_1;
    end
    if (_T_1) begin // @[yolo_layer.scala 430:50]
      temp2_index_0 <= 3'h0; // @[yolo_layer.scala 430:50]
    end else if (select2_0) begin // @[yolo_layer.scala 438:38]
      temp2_index_0 <= temp1_index_0;
    end else begin
      temp2_index_0 <= temp1_index_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  temp0_data_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  temp0_data_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  temp0_data_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  temp0_data_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  temp0_index_0 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  temp0_index_1 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  temp0_index_2 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  temp0_index_3 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  temp1_data_0 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  temp1_data_1 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  temp1_index_0 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  temp1_index_1 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  temp2_data_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  temp2_index_0 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module compare_2_cell(
  input         clock,
  input         reset,
  input  [31:0] io_data0,
  output [7:0]  io_max_data,
  output [6:0]  io_max_index
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] data0_cls_confidence = io_data0[7:0]; // @[yolo_layer.scala 370:40]
  wire [6:0] data0_cls_class = io_data0[14:8]; // @[yolo_layer.scala 371:35]
  reg [7:0] max_data; // @[yolo_layer.scala 375:27]
  reg [6:0] max_index; // @[yolo_layer.scala 376:28]
  wire  select = data0_cls_confidence > data0_cls_confidence; // @[yolo_layer.scala 381:40]
  assign io_max_data = max_data; // @[yolo_layer.scala 385:17]
  assign io_max_index = max_index; // @[yolo_layer.scala 386:18]
  always @(posedge clock) begin
    if (reset) begin // @[yolo_layer.scala 375:27]
      max_data <= 8'h0; // @[yolo_layer.scala 375:27]
    end else if (select) begin // @[yolo_layer.scala 383:20]
      max_data <= data0_cls_confidence;
    end else begin
      max_data <= data0_cls_confidence;
    end
    if (reset) begin // @[yolo_layer.scala 376:28]
      max_index <= 7'h0; // @[yolo_layer.scala 376:28]
    end else if (select) begin // @[yolo_layer.scala 384:21]
      max_index <= data0_cls_class;
    end else begin
      max_index <= data0_cls_class;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max_data = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  max_index = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module yolo_layer(
  input         clock,
  input         reset,
  input         io_yolo_layer_cls_en,
  output        io_yolo_cls_finish,
  input  [1:0]  io_yolo_current_cls_detect_layer,
  input  [3:0]  io_yolo_layer_cls_div_cnt,
  output [11:0] io_ofm_read_addr,
  input  [63:0] io_ofm_write_data_before,
  input         io_ofm_write_en_before,
  output [63:0] io_ofm_write_data_after,
  output        io_ofm_write_en_after,
  output [11:0] io_ofm_write_addr_after,
  output [7:0]  io_data_before_sigmoid,
  input  [23:0] io_data_after_sigmoid,
  output        io_sigmoid_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
`endif // RANDOMIZE_REG_INIT
  wire  unit_clock; // @[yolo_layer.scala 96:22]
  wire  unit_reset; // @[yolo_layer.scala 96:22]
  wire  unit_io_yolo_layer_finish; // @[yolo_layer.scala 96:22]
  wire [63:0] unit_io_data; // @[yolo_layer.scala 96:22]
  wire [7:0] unit_io_max_data; // @[yolo_layer.scala 96:22]
  wire [2:0] unit_io_max_index; // @[yolo_layer.scala 96:22]
  wire  cmp2_clock; // @[yolo_layer.scala 112:22]
  wire  cmp2_reset; // @[yolo_layer.scala 112:22]
  wire [31:0] cmp2_io_data0; // @[yolo_layer.scala 112:22]
  wire [7:0] cmp2_io_max_data; // @[yolo_layer.scala 112:22]
  wire [6:0] cmp2_io_max_index; // @[yolo_layer.scala 112:22]
  wire  yolo_layer_cls_last_div = io_yolo_layer_cls_div_cnt == 4'h9; // @[yolo_layer.scala 35:61]
  wire  sigmoid_en = yolo_layer_cls_last_div & io_yolo_layer_cls_en; // @[yolo_layer.scala 36:46]
  wire  cur_layer_sel_0 = io_yolo_current_cls_detect_layer == 2'h0; // @[yolo_layer.scala 39:103]
  wire  cur_layer_sel_1 = io_yolo_current_cls_detect_layer == 2'h1; // @[yolo_layer.scala 39:103]
  wire  cur_layer_sel_2 = io_yolo_current_cls_detect_layer == 2'h2; // @[yolo_layer.scala 39:103]
  wire [8:0] _anchor_number_T = cur_layer_sel_2 ? 9'h190 : 9'h0; // @[Mux.scala 101:16]
  wire [10:0] _anchor_number_T_1 = cur_layer_sel_1 ? 11'h640 : {{2'd0}, _anchor_number_T}; // @[Mux.scala 101:16]
  wire [12:0] anchor_number = cur_layer_sel_0 ? 13'h1900 : {{2'd0}, _anchor_number_T_1}; // @[Mux.scala 101:16]
  reg  ofm_write_data_sel_after_sigmoid_r_22; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_r; // @[Reg.scala 35:20]
  wire  ofm_write_data_sel_wire = sigmoid_en ? ofm_write_data_sel_after_sigmoid_r_22 : ofm_write_data_sel_r; // @[yolo_layer.scala 71:36]
  wire [12:0] _yolo_cls_finish_T_1 = anchor_number - 13'h1; // @[yolo_layer.scala 90:93]
  wire [12:0] _GEN_89 = {{1'd0}, io_ofm_write_addr_after}; // @[yolo_layer.scala 90:74]
  wire  _yolo_cls_finish_T_2 = _GEN_89 == _yolo_cls_finish_T_1; // @[yolo_layer.scala 90:74]
  wire  yolo_cls_finish = io_ofm_write_en_after & _GEN_89 == _yolo_cls_finish_T_1; // @[yolo_layer.scala 90:46]
  wire  _T_1 = reset | yolo_cls_finish; // @[yolo_layer.scala 76:28]
  reg [12:0] anchor_cnt_reg; // @[yolo_layer.scala 77:37]
  wire [12:0] _anchor_cnt_reg_T_5 = anchor_cnt_reg + 13'h1; // @[yolo_layer.scala 78:139]
  wire [11:0] ofm_read_addr = anchor_cnt_reg[12:1]; // @[yolo_layer.scala 82:32]
  reg [11:0] io_ofm_read_addr_r; // @[Reg.scala 35:20]
  reg [11:0] io_ofm_read_addr_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_r; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_r_2; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_r_3; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_r; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_r_1; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_r_2; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_r_3; // @[Reg.scala 35:20]
  wire  yolo_cls_part_finish = io_ofm_write_en_after & (io_ofm_write_addr_after == 12'he5f | _yolo_cls_finish_T_2); // @[yolo_layer.scala 88:51]
  wire  temp = anchor_cnt_reg[0]; // @[yolo_layer.scala 92:26]
  reg  ofm_read_data_sel_r; // @[Reg.scala 35:20]
  reg  ofm_read_data_sel_r_1; // @[Reg.scala 35:20]
  reg  ofm_read_data_sel_r_2; // @[Reg.scala 35:20]
  wire [6:0] _cls_part_max_index_entire_T = {io_yolo_layer_cls_div_cnt, 3'h0}; // @[yolo_layer.scala 107:83]
  wire [2:0] cls_part_max_index = unit_io_max_index; // @[yolo_layer.scala 101:24 44:34]
  wire [6:0] _GEN_91 = {{4'd0}, cls_part_max_index}; // @[yolo_layer.scala 107:54]
  wire [6:0] cls_part_max_index_entire = _GEN_91 + _cls_part_max_index_entire_T; // @[yolo_layer.scala 107:54]
  wire [23:0] data0_hi = {17'h0,cls_part_max_index_entire}; // @[Cat.scala 33:92]
  wire [7:0] cls_part_max_data = unit_io_max_data; // @[yolo_layer.scala 100:23 43:33]
  wire [6:0] max_index = cmp2_io_max_index; // @[yolo_layer.scala 111:25 117:15]
  wire [15:0] max_data_fp = io_data_after_sigmoid[15:0]; // @[yolo_layer.scala 121:27 122:17]
  wire [23:0] data_after_sigmoid = {1'h0,max_index,max_data_fp}; // @[Cat.scala 33:92]
  wire [7:0] max_data = cmp2_io_max_data; // @[yolo_layer.scala 110:24 116:14]
  wire [31:0] data_after_cmp2 = {17'h0,max_index,max_data}; // @[Cat.scala 33:92]
  wire  _ofm_after_cmp_data_0_T = ofm_write_en_after_r_3 & io_yolo_layer_cls_en; // @[yolo_layer.scala 131:89]
  reg [31:0] ofm_after_cmp_data_0_r; // @[Reg.scala 35:20]
  reg [31:0] ofm_after_cmp_data_1_r; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_22; // @[Reg.scala 35:20]
  reg [23:0] ofm_after_sigmoid_data_0_r; // @[Reg.scala 35:20]
  reg [31:0] ofm_after_sigmoid_data_1_r; // @[Reg.scala 35:20]
  wire [31:0] ofm_after_sigmoid_data_0 = {{8'd0}, ofm_after_sigmoid_data_0_r}; // @[yolo_layer.scala 127:38 139:39]
  wire [63:0] ofm_write_data_after_no_sigmoid = {ofm_after_cmp_data_1_r,ofm_after_cmp_data_0_r}; // @[Cat.scala 33:92]
  wire [63:0] ofm_write_data_after_has_sigmoid = {ofm_after_sigmoid_data_1_r,ofm_after_sigmoid_data_0}; // @[Cat.scala 33:92]
  reg  ofm_write_en_after_sigmoid_r; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_1; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_2; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_3; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_4; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_5; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_6; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_7; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_8; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_9; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_10; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_11; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_12; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_13; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_14; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_15; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_16; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_17; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_18; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_19; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_20; // @[Reg.scala 35:20]
  reg  ofm_write_en_after_sigmoid_r_21; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_1; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_2; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_3; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_4; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_5; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_6; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_7; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_8; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_9; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_10; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_11; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_12; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_13; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_14; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_15; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_16; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_17; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_18; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_19; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_20; // @[Reg.scala 35:20]
  reg  ofm_write_data_sel_after_sigmoid_r_21; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_1; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_2; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_3; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_4; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_5; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_6; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_7; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_8; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_9; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_10; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_11; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_12; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_13; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_14; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_15; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_16; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_17; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_18; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_19; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_20; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid_r_21; // @[Reg.scala 35:20]
  reg [11:0] ofm_write_addr_after_sigmoid; // @[Reg.scala 35:20]
  wire  ofm_write_en_after_wire = sigmoid_en ? ofm_write_en_after_sigmoid_r_22 : ofm_write_en_after_r_3; // @[yolo_layer.scala 155:38]
  reg [11:0] io_ofm_write_addr_after_REG; // @[yolo_layer.scala 160:37]
  reg  io_ofm_write_en_after_REG; // @[yolo_layer.scala 162:37]
  compare_8_cell unit ( // @[yolo_layer.scala 96:22]
    .clock(unit_clock),
    .reset(unit_reset),
    .io_yolo_layer_finish(unit_io_yolo_layer_finish),
    .io_data(unit_io_data),
    .io_max_data(unit_io_max_data),
    .io_max_index(unit_io_max_index)
  );
  compare_2_cell cmp2 ( // @[yolo_layer.scala 112:22]
    .clock(cmp2_clock),
    .reset(cmp2_reset),
    .io_data0(cmp2_io_data0),
    .io_max_data(cmp2_io_max_data),
    .io_max_index(cmp2_io_max_index)
  );
  assign io_yolo_cls_finish = cur_layer_sel_0 ? yolo_cls_part_finish : yolo_cls_finish; // @[yolo_layer.scala 87:30]
  assign io_ofm_read_addr = io_ofm_read_addr_r_1; // @[yolo_layer.scala 83:22]
  assign io_ofm_write_data_after = sigmoid_en ? ofm_write_data_after_has_sigmoid : ofm_write_data_after_no_sigmoid; // @[yolo_layer.scala 150:31]
  assign io_ofm_write_en_after = io_ofm_write_en_after_REG; // @[yolo_layer.scala 162:27]
  assign io_ofm_write_addr_after = io_ofm_write_addr_after_REG; // @[yolo_layer.scala 160:28]
  assign io_data_before_sigmoid = cmp2_io_max_data; // @[yolo_layer.scala 110:24 116:14]
  assign io_sigmoid_en = yolo_layer_cls_last_div & io_yolo_layer_cls_en; // @[yolo_layer.scala 36:46]
  assign unit_clock = clock;
  assign unit_reset = reset;
  assign unit_io_yolo_layer_finish = io_yolo_cls_finish; // @[yolo_layer.scala 98:31]
  assign unit_io_data = io_ofm_write_data_before; // @[yolo_layer.scala 99:18]
  assign cmp2_clock = clock;
  assign cmp2_reset = reset;
  assign cmp2_io_data0 = {data0_hi,cls_part_max_data}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_22 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_22 <= ofm_write_data_sel_after_sigmoid_r_21; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_r <= ofm_read_data_sel_r_2; // @[Reg.scala 36:22]
    end
    if (_T_1) begin // @[yolo_layer.scala 77:37]
      anchor_cnt_reg <= 13'h0; // @[yolo_layer.scala 77:37]
    end else if (io_ofm_write_en_before & io_yolo_layer_cls_en) begin // @[yolo_layer.scala 78:30]
      if (anchor_cnt_reg != _yolo_cls_finish_T_1) begin // @[yolo_layer.scala 78:81]
        anchor_cnt_reg <= _anchor_cnt_reg_T_5;
      end else begin
        anchor_cnt_reg <= 13'h0;
      end
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_ofm_read_addr_r <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      io_ofm_read_addr_r <= ofm_read_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      io_ofm_read_addr_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      io_ofm_read_addr_r_1 <= io_ofm_read_addr_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_r <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_r <= ofm_read_addr; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_r_1 <= ofm_write_addr_after_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_r_2 <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_r_2 <= ofm_write_addr_after_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_r_3 <= 12'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_r_3 <= ofm_write_addr_after_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_r <= io_ofm_write_en_before; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_r_1 <= ofm_write_en_after_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_r_2 <= ofm_write_en_after_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_r_3 <= ofm_write_en_after_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_read_data_sel_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_read_data_sel_r <= temp; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_read_data_sel_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_read_data_sel_r_1 <= ofm_read_data_sel_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_read_data_sel_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else if (io_yolo_layer_cls_en) begin // @[Reg.scala 36:18]
      ofm_read_data_sel_r_2 <= ofm_read_data_sel_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_after_cmp_data_0_r <= 32'h0; // @[Reg.scala 35:20]
    end else if (_ofm_after_cmp_data_0_T) begin // @[Reg.scala 36:18]
      ofm_after_cmp_data_0_r <= data_after_cmp2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_after_cmp_data_1_r <= 32'h0; // @[Reg.scala 35:20]
    end else if (_ofm_after_cmp_data_0_T) begin // @[Reg.scala 36:18]
      ofm_after_cmp_data_1_r <= ofm_after_cmp_data_0_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_22 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_22 <= ofm_write_en_after_sigmoid_r_21; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_after_sigmoid_data_0_r <= 24'h0; // @[Reg.scala 35:20]
    end else if (ofm_write_en_after_sigmoid_r_22) begin // @[Reg.scala 36:18]
      ofm_after_sigmoid_data_0_r <= data_after_sigmoid; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_after_sigmoid_data_1_r <= 32'h0; // @[Reg.scala 35:20]
    end else if (ofm_write_en_after_sigmoid_r_22) begin // @[Reg.scala 36:18]
      ofm_after_sigmoid_data_1_r <= ofm_after_sigmoid_data_0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r <= ofm_write_en_after_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_1 <= ofm_write_en_after_sigmoid_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_2 <= ofm_write_en_after_sigmoid_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_3 <= ofm_write_en_after_sigmoid_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_4 <= ofm_write_en_after_sigmoid_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_5 <= ofm_write_en_after_sigmoid_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_6 <= ofm_write_en_after_sigmoid_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_7 <= ofm_write_en_after_sigmoid_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_8 <= ofm_write_en_after_sigmoid_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_9 <= ofm_write_en_after_sigmoid_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_10 <= ofm_write_en_after_sigmoid_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_11 <= ofm_write_en_after_sigmoid_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_12 <= ofm_write_en_after_sigmoid_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_13 <= ofm_write_en_after_sigmoid_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_14 <= ofm_write_en_after_sigmoid_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_15 <= ofm_write_en_after_sigmoid_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_16 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_16 <= ofm_write_en_after_sigmoid_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_17 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_17 <= ofm_write_en_after_sigmoid_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_18 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_18 <= ofm_write_en_after_sigmoid_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_19 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_19 <= ofm_write_en_after_sigmoid_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_20 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_20 <= ofm_write_en_after_sigmoid_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_en_after_sigmoid_r_21 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_en_after_sigmoid_r_21 <= ofm_write_en_after_sigmoid_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r <= ofm_write_data_sel_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_1 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_1 <= ofm_write_data_sel_after_sigmoid_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_2 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_2 <= ofm_write_data_sel_after_sigmoid_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_3 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_3 <= ofm_write_data_sel_after_sigmoid_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_4 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_4 <= ofm_write_data_sel_after_sigmoid_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_5 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_5 <= ofm_write_data_sel_after_sigmoid_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_6 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_6 <= ofm_write_data_sel_after_sigmoid_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_7 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_7 <= ofm_write_data_sel_after_sigmoid_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_8 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_8 <= ofm_write_data_sel_after_sigmoid_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_9 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_9 <= ofm_write_data_sel_after_sigmoid_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_10 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_10 <= ofm_write_data_sel_after_sigmoid_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_11 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_11 <= ofm_write_data_sel_after_sigmoid_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_12 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_12 <= ofm_write_data_sel_after_sigmoid_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_13 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_13 <= ofm_write_data_sel_after_sigmoid_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_14 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_14 <= ofm_write_data_sel_after_sigmoid_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_15 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_15 <= ofm_write_data_sel_after_sigmoid_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_16 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_16 <= ofm_write_data_sel_after_sigmoid_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_17 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_17 <= ofm_write_data_sel_after_sigmoid_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_18 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_18 <= ofm_write_data_sel_after_sigmoid_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_19 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_19 <= ofm_write_data_sel_after_sigmoid_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_20 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_20 <= ofm_write_data_sel_after_sigmoid_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_data_sel_after_sigmoid_r_21 <= 1'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_data_sel_after_sigmoid_r_21 <= ofm_write_data_sel_after_sigmoid_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r <= ofm_write_addr_after_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_1 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_1 <= ofm_write_addr_after_sigmoid_r; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_2 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_2 <= ofm_write_addr_after_sigmoid_r_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_3 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_3 <= ofm_write_addr_after_sigmoid_r_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_4 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_4 <= ofm_write_addr_after_sigmoid_r_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_5 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_5 <= ofm_write_addr_after_sigmoid_r_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_6 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_6 <= ofm_write_addr_after_sigmoid_r_5; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_7 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_7 <= ofm_write_addr_after_sigmoid_r_6; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_8 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_8 <= ofm_write_addr_after_sigmoid_r_7; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_9 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_9 <= ofm_write_addr_after_sigmoid_r_8; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_10 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_10 <= ofm_write_addr_after_sigmoid_r_9; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_11 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_11 <= ofm_write_addr_after_sigmoid_r_10; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_12 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_12 <= ofm_write_addr_after_sigmoid_r_11; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_13 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_13 <= ofm_write_addr_after_sigmoid_r_12; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_14 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_14 <= ofm_write_addr_after_sigmoid_r_13; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_15 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_15 <= ofm_write_addr_after_sigmoid_r_14; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_16 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_16 <= ofm_write_addr_after_sigmoid_r_15; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_17 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_17 <= ofm_write_addr_after_sigmoid_r_16; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_18 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_18 <= ofm_write_addr_after_sigmoid_r_17; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_19 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_19 <= ofm_write_addr_after_sigmoid_r_18; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_20 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_20 <= ofm_write_addr_after_sigmoid_r_19; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid_r_21 <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid_r_21 <= ofm_write_addr_after_sigmoid_r_20; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      ofm_write_addr_after_sigmoid <= 12'h0; // @[Reg.scala 35:20]
    end else if (sigmoid_en) begin // @[Reg.scala 36:18]
      ofm_write_addr_after_sigmoid <= ofm_write_addr_after_sigmoid_r_21; // @[Reg.scala 36:22]
    end
    if (sigmoid_en) begin // @[yolo_layer.scala 160:41]
      io_ofm_write_addr_after_REG <= ofm_write_addr_after_sigmoid;
    end else begin
      io_ofm_write_addr_after_REG <= ofm_write_addr_after_r_3;
    end
    io_ofm_write_en_after_REG <= ofm_write_en_after_wire & ofm_write_data_sel_wire; // @[yolo_layer.scala 162:62]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_22 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ofm_write_data_sel_r = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  anchor_cnt_reg = _RAND_2[12:0];
  _RAND_3 = {1{`RANDOM}};
  io_ofm_read_addr_r = _RAND_3[11:0];
  _RAND_4 = {1{`RANDOM}};
  io_ofm_read_addr_r_1 = _RAND_4[11:0];
  _RAND_5 = {1{`RANDOM}};
  ofm_write_addr_after_r = _RAND_5[11:0];
  _RAND_6 = {1{`RANDOM}};
  ofm_write_addr_after_r_1 = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  ofm_write_addr_after_r_2 = _RAND_7[11:0];
  _RAND_8 = {1{`RANDOM}};
  ofm_write_addr_after_r_3 = _RAND_8[11:0];
  _RAND_9 = {1{`RANDOM}};
  ofm_write_en_after_r = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ofm_write_en_after_r_1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ofm_write_en_after_r_2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ofm_write_en_after_r_3 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ofm_read_data_sel_r = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  ofm_read_data_sel_r_1 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  ofm_read_data_sel_r_2 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  ofm_after_cmp_data_0_r = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  ofm_after_cmp_data_1_r = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_22 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ofm_after_sigmoid_data_0_r = _RAND_19[23:0];
  _RAND_20 = {1{`RANDOM}};
  ofm_after_sigmoid_data_1_r = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_5 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_6 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_7 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_8 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_9 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_10 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_11 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_12 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_13 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_14 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_15 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_16 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_17 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_18 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_19 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_20 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  ofm_write_en_after_sigmoid_r_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_1 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_2 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_3 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_4 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_5 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_6 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_7 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_8 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_9 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_10 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_11 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_12 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_13 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_14 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_15 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_16 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_17 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_18 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_19 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_20 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  ofm_write_data_sel_after_sigmoid_r_21 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r = _RAND_65[11:0];
  _RAND_66 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_1 = _RAND_66[11:0];
  _RAND_67 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_2 = _RAND_67[11:0];
  _RAND_68 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_3 = _RAND_68[11:0];
  _RAND_69 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_4 = _RAND_69[11:0];
  _RAND_70 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_5 = _RAND_70[11:0];
  _RAND_71 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_6 = _RAND_71[11:0];
  _RAND_72 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_7 = _RAND_72[11:0];
  _RAND_73 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_8 = _RAND_73[11:0];
  _RAND_74 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_9 = _RAND_74[11:0];
  _RAND_75 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_10 = _RAND_75[11:0];
  _RAND_76 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_11 = _RAND_76[11:0];
  _RAND_77 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_12 = _RAND_77[11:0];
  _RAND_78 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_13 = _RAND_78[11:0];
  _RAND_79 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_14 = _RAND_79[11:0];
  _RAND_80 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_15 = _RAND_80[11:0];
  _RAND_81 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_16 = _RAND_81[11:0];
  _RAND_82 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_17 = _RAND_82[11:0];
  _RAND_83 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_18 = _RAND_83[11:0];
  _RAND_84 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_19 = _RAND_84[11:0];
  _RAND_85 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_20 = _RAND_85[11:0];
  _RAND_86 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid_r_21 = _RAND_86[11:0];
  _RAND_87 = {1{`RANDOM}};
  ofm_write_addr_after_sigmoid = _RAND_87[11:0];
  _RAND_88 = {1{`RANDOM}};
  io_ofm_write_addr_after_REG = _RAND_88[11:0];
  _RAND_89 = {1{`RANDOM}};
  io_ofm_write_en_after_REG = _RAND_89[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module sint2float(
  input         clock,
  input         reset,
  input         io_i_valid,
  input  [31:0] io_i_data,
  output [31:0] io_o_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  i_sign; // @[Arithmetic.scala 26:23]
  reg [30:0] i_uint; // @[Arithmetic.scala 27:23]
  wire [30:0] _i_uint_T_2 = ~io_i_data[30:0]; // @[Arithmetic.scala 30:35]
  wire [30:0] _i_uint_T_4 = _i_uint_T_2 + 31'h1; // @[Arithmetic.scala 30:61]
  reg  float_sign; // @[Arithmetic.scala 33:27]
  reg [7:0] float_exp; // @[Arithmetic.scala 34:27]
  reg [22:0] float_frac; // @[Arithmetic.scala 35:27]
  reg  REG; // @[Arithmetic.scala 36:15]
  wire [53:0] data_extend = {i_uint,23'h0}; // @[Cat.scala 33:92]
  wire [22:0] _GEN_2 = i_uint[0] ? data_extend[22:0] : 23'h0; // @[Arithmetic.scala 39:16 42:30 43:20]
  wire [6:0] _GEN_3 = i_uint[0] ? 7'h7f : 7'h0; // @[Arithmetic.scala 38:16 42:30 44:20]
  wire [22:0] _GEN_4 = i_uint[1] ? data_extend[23:1] : _GEN_2; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_5 = i_uint[1] ? 8'h80 : {{1'd0}, _GEN_3}; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_6 = i_uint[2] ? data_extend[24:2] : _GEN_4; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_7 = i_uint[2] ? 8'h81 : _GEN_5; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_8 = i_uint[3] ? data_extend[25:3] : _GEN_6; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_9 = i_uint[3] ? 8'h82 : _GEN_7; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_10 = i_uint[4] ? data_extend[26:4] : _GEN_8; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_11 = i_uint[4] ? 8'h83 : _GEN_9; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_12 = i_uint[5] ? data_extend[27:5] : _GEN_10; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_13 = i_uint[5] ? 8'h84 : _GEN_11; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_14 = i_uint[6] ? data_extend[28:6] : _GEN_12; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_15 = i_uint[6] ? 8'h85 : _GEN_13; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_16 = i_uint[7] ? data_extend[29:7] : _GEN_14; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_17 = i_uint[7] ? 8'h86 : _GEN_15; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_18 = i_uint[8] ? data_extend[30:8] : _GEN_16; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_19 = i_uint[8] ? 8'h87 : _GEN_17; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_20 = i_uint[9] ? data_extend[31:9] : _GEN_18; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_21 = i_uint[9] ? 8'h88 : _GEN_19; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_22 = i_uint[10] ? data_extend[32:10] : _GEN_20; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_23 = i_uint[10] ? 8'h89 : _GEN_21; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_24 = i_uint[11] ? data_extend[33:11] : _GEN_22; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_25 = i_uint[11] ? 8'h8a : _GEN_23; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_26 = i_uint[12] ? data_extend[34:12] : _GEN_24; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_27 = i_uint[12] ? 8'h8b : _GEN_25; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_28 = i_uint[13] ? data_extend[35:13] : _GEN_26; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_29 = i_uint[13] ? 8'h8c : _GEN_27; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_30 = i_uint[14] ? data_extend[36:14] : _GEN_28; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_31 = i_uint[14] ? 8'h8d : _GEN_29; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_32 = i_uint[15] ? data_extend[37:15] : _GEN_30; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_33 = i_uint[15] ? 8'h8e : _GEN_31; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_34 = i_uint[16] ? data_extend[38:16] : _GEN_32; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_35 = i_uint[16] ? 8'h8f : _GEN_33; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_36 = i_uint[17] ? data_extend[39:17] : _GEN_34; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_37 = i_uint[17] ? 8'h90 : _GEN_35; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_38 = i_uint[18] ? data_extend[40:18] : _GEN_36; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_39 = i_uint[18] ? 8'h91 : _GEN_37; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_40 = i_uint[19] ? data_extend[41:19] : _GEN_38; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_41 = i_uint[19] ? 8'h92 : _GEN_39; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_42 = i_uint[20] ? data_extend[42:20] : _GEN_40; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_43 = i_uint[20] ? 8'h93 : _GEN_41; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_44 = i_uint[21] ? data_extend[43:21] : _GEN_42; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_45 = i_uint[21] ? 8'h94 : _GEN_43; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_46 = i_uint[22] ? data_extend[44:22] : _GEN_44; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_47 = i_uint[22] ? 8'h95 : _GEN_45; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_48 = i_uint[23] ? data_extend[45:23] : _GEN_46; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_49 = i_uint[23] ? 8'h96 : _GEN_47; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_50 = i_uint[24] ? data_extend[46:24] : _GEN_48; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_51 = i_uint[24] ? 8'h97 : _GEN_49; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_52 = i_uint[25] ? data_extend[47:25] : _GEN_50; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_53 = i_uint[25] ? 8'h98 : _GEN_51; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_54 = i_uint[26] ? data_extend[48:26] : _GEN_52; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_55 = i_uint[26] ? 8'h99 : _GEN_53; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_56 = i_uint[27] ? data_extend[49:27] : _GEN_54; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_57 = i_uint[27] ? 8'h9a : _GEN_55; // @[Arithmetic.scala 42:30 44:20]
  wire [22:0] _GEN_58 = i_uint[28] ? data_extend[50:28] : _GEN_56; // @[Arithmetic.scala 42:30 43:20]
  wire [7:0] _GEN_59 = i_uint[28] ? 8'h9b : _GEN_57; // @[Arithmetic.scala 42:30 44:20]
  wire [8:0] io_o_data_hi = {float_sign,float_exp}; // @[Cat.scala 33:92]
  assign io_o_data = {io_o_data_hi,float_frac}; // @[Cat.scala 33:92]
  always @(posedge clock) begin
    if (reset) begin // @[Arithmetic.scala 26:23]
      i_sign <= 1'h0; // @[Arithmetic.scala 26:23]
    end else if (io_i_valid) begin // @[Arithmetic.scala 28:20]
      i_sign <= io_i_data[31]; // @[Arithmetic.scala 29:12]
    end
    if (reset) begin // @[Arithmetic.scala 27:23]
      i_uint <= 31'h0; // @[Arithmetic.scala 27:23]
    end else if (io_i_valid) begin // @[Arithmetic.scala 28:20]
      if (io_i_data[31]) begin // @[Arithmetic.scala 30:18]
        i_uint <= _i_uint_T_4;
      end else begin
        i_uint <= io_i_data[30:0];
      end
    end
    if (reset) begin // @[Arithmetic.scala 33:27]
      float_sign <= 1'h0; // @[Arithmetic.scala 33:27]
    end else if (REG) begin // @[Arithmetic.scala 36:32]
      float_sign <= i_sign; // @[Arithmetic.scala 37:16]
    end
    if (reset) begin // @[Arithmetic.scala 34:27]
      float_exp <= 8'h0; // @[Arithmetic.scala 34:27]
    end else if (REG) begin // @[Arithmetic.scala 36:32]
      if (i_uint[30]) begin // @[Arithmetic.scala 42:30]
        float_exp <= 8'h9d; // @[Arithmetic.scala 44:20]
      end else if (i_uint[29]) begin // @[Arithmetic.scala 42:30]
        float_exp <= 8'h9c; // @[Arithmetic.scala 44:20]
      end else begin
        float_exp <= _GEN_59;
      end
    end
    if (reset) begin // @[Arithmetic.scala 35:27]
      float_frac <= 23'h0; // @[Arithmetic.scala 35:27]
    end else if (REG) begin // @[Arithmetic.scala 36:32]
      if (i_uint[30]) begin // @[Arithmetic.scala 42:30]
        float_frac <= data_extend[52:30]; // @[Arithmetic.scala 43:20]
      end else if (i_uint[29]) begin // @[Arithmetic.scala 42:30]
        float_frac <= data_extend[51:29]; // @[Arithmetic.scala 43:20]
      end else begin
        float_frac <= _GEN_58;
      end
    end
    if (reset) begin // @[Arithmetic.scala 36:15]
      REG <= 1'h0; // @[Arithmetic.scala 36:15]
    end else begin
      REG <= io_i_valid; // @[Arithmetic.scala 36:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_sign = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  i_uint = _RAND_1[30:0];
  _RAND_2 = {1{`RANDOM}};
  float_sign = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  float_exp = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  float_frac = _RAND_4[22:0];
  _RAND_5 = {1{`RANDOM}};
  REG = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP32_Mult(
  input         clock,
  input         reset,
  input  [31:0] io_x,
  input  [31:0] io_y,
  output [31:0] io_z,
  input         io_valid_in
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  zs = io_x[31] ^ io_y[31]; // @[FP32.scala 179:21]
  wire [7:0] xe = io_x[30:23]; // @[FP32.scala 180:16]
  wire [7:0] ye = io_y[30:23]; // @[FP32.scala 181:16]
  wire [22:0] xf = io_x[22:0]; // @[FP32.scala 182:16]
  wire [22:0] yf = io_y[22:0]; // @[FP32.scala 183:16]
  wire  _is_zero_T_2 = xe == 8'h0 | ye == 8'h0; // @[FP32.scala 185:38]
  reg  is_zero; // @[Reg.scala 19:16]
  wire [23:0] _zf_0_T = {1'h1,xf}; // @[Cat.scala 33:92]
  wire [23:0] _zf_0_T_1 = {1'h1,yf}; // @[Cat.scala 33:92]
  wire [47:0] _zf_0_T_2 = _zf_0_T * _zf_0_T_1; // @[FP32.scala 187:28]
  wire [25:0] zf_0 = _zf_0_T_2[47:22]; // @[FP32.scala 187:43]
  reg [24:0] zf_1; // @[Reg.scala 19:16]
  reg  valid_in_r; // @[FP32.scala 190:27]
  reg  carry_r; // @[Reg.scala 19:16]
  wire  carry = carry_r | zf_1 == 25'h1ffffff; // @[FP32.scala 192:48]
  wire [22:0] _GEN_6 = {{22'd0}, zf_1[1]}; // @[FP32.scala 193:38]
  wire [22:0] _zf_T_3 = zf_1[24:2] + _GEN_6; // @[FP32.scala 193:38]
  wire [22:0] _GEN_7 = {{22'd0}, zf_1[0]}; // @[FP32.scala 193:61]
  wire [22:0] _zf_T_7 = zf_1[23:1] + _GEN_7; // @[FP32.scala 193:61]
  wire [22:0] zf = carry ? _zf_T_3 : _zf_T_7; // @[FP32.scala 193:18]
  wire [7:0] _ze_T_1 = xe + ye; // @[FP32.scala 194:28]
  reg [7:0] ze_r; // @[Reg.scala 19:16]
  wire [6:0] _ze_T_2 = carry ? 7'h7e : 7'h7f; // @[FP32.scala 194:52]
  wire [7:0] _GEN_8 = {{1'd0}, _ze_T_2}; // @[FP32.scala 194:47]
  wire [7:0] ze = ze_r - _GEN_8; // @[FP32.scala 194:47]
  reg  out_z_r; // @[Reg.scala 19:16]
  wire [30:0] _out_z_T_1 = {ze,zf}; // @[Cat.scala 33:92]
  wire [30:0] _out_z_T_2 = is_zero ? 31'h0 : _out_z_T_1; // @[Mux.scala 47:70]
  wire [31:0] out_z = {out_z_r,_out_z_T_2}; // @[Cat.scala 33:92]
  reg [31:0] io_z_r; // @[Reg.scala 19:16]
  assign io_z = io_z_r; // @[FP32.scala 207:8]
  always @(posedge clock) begin
    if (io_valid_in) begin // @[Reg.scala 20:18]
      is_zero <= _is_zero_T_2; // @[Reg.scala 20:22]
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      zf_1 <= zf_0[24:0]; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[FP32.scala 190:27]
      valid_in_r <= 1'h0; // @[FP32.scala 190:27]
    end else begin
      valid_in_r <= io_valid_in; // @[FP32.scala 190:27]
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      carry_r <= zf_0[25]; // @[Reg.scala 20:22]
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      ze_r <= _ze_T_1; // @[Reg.scala 20:22]
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      out_z_r <= zs; // @[Reg.scala 20:22]
    end
    if (valid_in_r) begin // @[Reg.scala 20:18]
      io_z_r <= out_z; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  is_zero = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  zf_1 = _RAND_1[24:0];
  _RAND_2 = {1{`RANDOM}};
  valid_in_r = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  carry_r = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ze_r = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  out_z_r = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  io_z_r = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dequant_cell(
  input         clock,
  input         reset,
  input         io_en,
  input  [7:0]  io_i_data,
  input  [31:0] io_scale,
  output [31:0] io_o_data,
  input  [7:0]  io_zero_point
);
  wire  sub_module_clock; // @[act.scala 221:28]
  wire  sub_module_reset; // @[act.scala 221:28]
  wire [7:0] sub_module_io_zero_point; // @[act.scala 221:28]
  wire [7:0] sub_module_io_data_in; // @[act.scala 221:28]
  wire [7:0] sub_module_io_data_out; // @[act.scala 221:28]
  wire  convert_data_convert_clock; // @[Arithmetic.scala 77:27]
  wire  convert_data_convert_reset; // @[Arithmetic.scala 77:27]
  wire  convert_data_convert_io_i_valid; // @[Arithmetic.scala 77:27]
  wire [31:0] convert_data_convert_io_i_data; // @[Arithmetic.scala 77:27]
  wire [31:0] convert_data_convert_io_o_data; // @[Arithmetic.scala 77:27]
  wire  fp32_data_muler_clock; // @[Arithmetic.scala 95:25]
  wire  fp32_data_muler_reset; // @[Arithmetic.scala 95:25]
  wire [31:0] fp32_data_muler_io_x; // @[Arithmetic.scala 95:25]
  wire [31:0] fp32_data_muler_io_y; // @[Arithmetic.scala 95:25]
  wire [31:0] fp32_data_muler_io_z; // @[Arithmetic.scala 95:25]
  wire  fp32_data_muler_io_valid_in; // @[Arithmetic.scala 95:25]
  wire [7:0] sub_out = sub_module_io_data_out; // @[act.scala 220:23 224:13]
  wire [23:0] _i_data_T_2 = sub_out[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 77:12]
  cal_sub_zero_point sub_module ( // @[act.scala 221:28]
    .clock(sub_module_clock),
    .reset(sub_module_reset),
    .io_zero_point(sub_module_io_zero_point),
    .io_data_in(sub_module_io_data_in),
    .io_data_out(sub_module_io_data_out)
  );
  sint2float convert_data_convert ( // @[Arithmetic.scala 77:27]
    .clock(convert_data_convert_clock),
    .reset(convert_data_convert_reset),
    .io_i_valid(convert_data_convert_io_i_valid),
    .io_i_data(convert_data_convert_io_i_data),
    .io_o_data(convert_data_convert_io_o_data)
  );
  FP32_Mult fp32_data_muler ( // @[Arithmetic.scala 95:25]
    .clock(fp32_data_muler_clock),
    .reset(fp32_data_muler_reset),
    .io_x(fp32_data_muler_io_x),
    .io_y(fp32_data_muler_io_y),
    .io_z(fp32_data_muler_io_z),
    .io_valid_in(fp32_data_muler_io_valid_in)
  );
  assign io_o_data = fp32_data_muler_io_z; // @[Arithmetic.scala 124:22 125:17]
  assign sub_module_clock = clock;
  assign sub_module_reset = reset;
  assign sub_module_io_zero_point = io_zero_point; // @[act.scala 222:30]
  assign sub_module_io_data_in = io_i_data; // @[act.scala 223:27]
  assign convert_data_convert_clock = clock;
  assign convert_data_convert_reset = reset;
  assign convert_data_convert_io_i_valid = io_en; // @[Arithmetic.scala 79:28]
  assign convert_data_convert_io_i_data = {_i_data_T_2,sub_out}; // @[Arithmetic.scala 78:30]
  assign fp32_data_muler_clock = clock;
  assign fp32_data_muler_reset = reset;
  assign fp32_data_muler_io_x = convert_data_convert_io_o_data; // @[Arithmetic.scala 124:22 125:17]
  assign fp32_data_muler_io_y = io_scale; // @[Arithmetic.scala 124:22 125:17]
  assign fp32_data_muler_io_valid_in = io_en; // @[Arithmetic.scala 98:25]
endmodule
module dequant_int8_2_fp32(
  input         clock,
  input         reset,
  input         io_en,
  input  [7:0]  io_i_data_0,
  input  [7:0]  io_i_data_1,
  input  [7:0]  io_i_data_2,
  input  [7:0]  io_i_data_3,
  input  [7:0]  io_i_data_4,
  input  [7:0]  io_i_data_5,
  input  [7:0]  io_i_data_6,
  input  [7:0]  io_i_data_7,
  input  [31:0] io_scale,
  input  [7:0]  io_zero_point,
  output [31:0] io_o_data_0,
  output [31:0] io_o_data_1,
  output [31:0] io_o_data_2,
  output [31:0] io_o_data_3,
  output [31:0] io_o_data_4,
  output [31:0] io_o_data_5,
  output [31:0] io_o_data_6,
  output [31:0] io_o_data_7
);
  wire  cell_0_clock; // @[act.scala 60:36]
  wire  cell_0_reset; // @[act.scala 60:36]
  wire  cell_0_io_en; // @[act.scala 60:36]
  wire [7:0] cell_0_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_0_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_0_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_0_io_zero_point; // @[act.scala 60:36]
  wire  cell_1_clock; // @[act.scala 60:36]
  wire  cell_1_reset; // @[act.scala 60:36]
  wire  cell_1_io_en; // @[act.scala 60:36]
  wire [7:0] cell_1_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_1_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_1_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_1_io_zero_point; // @[act.scala 60:36]
  wire  cell_2_clock; // @[act.scala 60:36]
  wire  cell_2_reset; // @[act.scala 60:36]
  wire  cell_2_io_en; // @[act.scala 60:36]
  wire [7:0] cell_2_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_2_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_2_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_2_io_zero_point; // @[act.scala 60:36]
  wire  cell_3_clock; // @[act.scala 60:36]
  wire  cell_3_reset; // @[act.scala 60:36]
  wire  cell_3_io_en; // @[act.scala 60:36]
  wire [7:0] cell_3_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_3_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_3_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_3_io_zero_point; // @[act.scala 60:36]
  wire  cell_4_clock; // @[act.scala 60:36]
  wire  cell_4_reset; // @[act.scala 60:36]
  wire  cell_4_io_en; // @[act.scala 60:36]
  wire [7:0] cell_4_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_4_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_4_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_4_io_zero_point; // @[act.scala 60:36]
  wire  cell_5_clock; // @[act.scala 60:36]
  wire  cell_5_reset; // @[act.scala 60:36]
  wire  cell_5_io_en; // @[act.scala 60:36]
  wire [7:0] cell_5_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_5_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_5_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_5_io_zero_point; // @[act.scala 60:36]
  wire  cell_6_clock; // @[act.scala 60:36]
  wire  cell_6_reset; // @[act.scala 60:36]
  wire  cell_6_io_en; // @[act.scala 60:36]
  wire [7:0] cell_6_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_6_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_6_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_6_io_zero_point; // @[act.scala 60:36]
  wire  cell_7_clock; // @[act.scala 60:36]
  wire  cell_7_reset; // @[act.scala 60:36]
  wire  cell_7_io_en; // @[act.scala 60:36]
  wire [7:0] cell_7_io_i_data; // @[act.scala 60:36]
  wire [31:0] cell_7_io_scale; // @[act.scala 60:36]
  wire [31:0] cell_7_io_o_data; // @[act.scala 60:36]
  wire [7:0] cell_7_io_zero_point; // @[act.scala 60:36]
  dequant_cell cell_0 ( // @[act.scala 60:36]
    .clock(cell_0_clock),
    .reset(cell_0_reset),
    .io_en(cell_0_io_en),
    .io_i_data(cell_0_io_i_data),
    .io_scale(cell_0_io_scale),
    .io_o_data(cell_0_io_o_data),
    .io_zero_point(cell_0_io_zero_point)
  );
  dequant_cell cell_1 ( // @[act.scala 60:36]
    .clock(cell_1_clock),
    .reset(cell_1_reset),
    .io_en(cell_1_io_en),
    .io_i_data(cell_1_io_i_data),
    .io_scale(cell_1_io_scale),
    .io_o_data(cell_1_io_o_data),
    .io_zero_point(cell_1_io_zero_point)
  );
  dequant_cell cell_2 ( // @[act.scala 60:36]
    .clock(cell_2_clock),
    .reset(cell_2_reset),
    .io_en(cell_2_io_en),
    .io_i_data(cell_2_io_i_data),
    .io_scale(cell_2_io_scale),
    .io_o_data(cell_2_io_o_data),
    .io_zero_point(cell_2_io_zero_point)
  );
  dequant_cell cell_3 ( // @[act.scala 60:36]
    .clock(cell_3_clock),
    .reset(cell_3_reset),
    .io_en(cell_3_io_en),
    .io_i_data(cell_3_io_i_data),
    .io_scale(cell_3_io_scale),
    .io_o_data(cell_3_io_o_data),
    .io_zero_point(cell_3_io_zero_point)
  );
  dequant_cell cell_4 ( // @[act.scala 60:36]
    .clock(cell_4_clock),
    .reset(cell_4_reset),
    .io_en(cell_4_io_en),
    .io_i_data(cell_4_io_i_data),
    .io_scale(cell_4_io_scale),
    .io_o_data(cell_4_io_o_data),
    .io_zero_point(cell_4_io_zero_point)
  );
  dequant_cell cell_5 ( // @[act.scala 60:36]
    .clock(cell_5_clock),
    .reset(cell_5_reset),
    .io_en(cell_5_io_en),
    .io_i_data(cell_5_io_i_data),
    .io_scale(cell_5_io_scale),
    .io_o_data(cell_5_io_o_data),
    .io_zero_point(cell_5_io_zero_point)
  );
  dequant_cell cell_6 ( // @[act.scala 60:36]
    .clock(cell_6_clock),
    .reset(cell_6_reset),
    .io_en(cell_6_io_en),
    .io_i_data(cell_6_io_i_data),
    .io_scale(cell_6_io_scale),
    .io_o_data(cell_6_io_o_data),
    .io_zero_point(cell_6_io_zero_point)
  );
  dequant_cell cell_7 ( // @[act.scala 60:36]
    .clock(cell_7_clock),
    .reset(cell_7_reset),
    .io_en(cell_7_io_en),
    .io_i_data(cell_7_io_i_data),
    .io_scale(cell_7_io_scale),
    .io_o_data(cell_7_io_o_data),
    .io_zero_point(cell_7_io_zero_point)
  );
  assign io_o_data_0 = cell_0_io_o_data; // @[act.scala 66:21]
  assign io_o_data_1 = cell_1_io_o_data; // @[act.scala 66:21]
  assign io_o_data_2 = cell_2_io_o_data; // @[act.scala 66:21]
  assign io_o_data_3 = cell_3_io_o_data; // @[act.scala 66:21]
  assign io_o_data_4 = cell_4_io_o_data; // @[act.scala 66:21]
  assign io_o_data_5 = cell_5_io_o_data; // @[act.scala 66:21]
  assign io_o_data_6 = cell_6_io_o_data; // @[act.scala 66:21]
  assign io_o_data_7 = cell_7_io_o_data; // @[act.scala 66:21]
  assign cell_0_clock = clock;
  assign cell_0_reset = reset;
  assign cell_0_io_en = io_en; // @[act.scala 62:22]
  assign cell_0_io_i_data = io_i_data_0; // @[act.scala 63:26]
  assign cell_0_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_0_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_1_clock = clock;
  assign cell_1_reset = reset;
  assign cell_1_io_en = io_en; // @[act.scala 62:22]
  assign cell_1_io_i_data = io_i_data_1; // @[act.scala 63:26]
  assign cell_1_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_1_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_2_clock = clock;
  assign cell_2_reset = reset;
  assign cell_2_io_en = io_en; // @[act.scala 62:22]
  assign cell_2_io_i_data = io_i_data_2; // @[act.scala 63:26]
  assign cell_2_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_2_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_3_clock = clock;
  assign cell_3_reset = reset;
  assign cell_3_io_en = io_en; // @[act.scala 62:22]
  assign cell_3_io_i_data = io_i_data_3; // @[act.scala 63:26]
  assign cell_3_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_3_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_4_clock = clock;
  assign cell_4_reset = reset;
  assign cell_4_io_en = io_en; // @[act.scala 62:22]
  assign cell_4_io_i_data = io_i_data_4; // @[act.scala 63:26]
  assign cell_4_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_4_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_5_clock = clock;
  assign cell_5_reset = reset;
  assign cell_5_io_en = io_en; // @[act.scala 62:22]
  assign cell_5_io_i_data = io_i_data_5; // @[act.scala 63:26]
  assign cell_5_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_5_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_6_clock = clock;
  assign cell_6_reset = reset;
  assign cell_6_io_en = io_en; // @[act.scala 62:22]
  assign cell_6_io_i_data = io_i_data_6; // @[act.scala 63:26]
  assign cell_6_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_6_io_zero_point = io_zero_point; // @[act.scala 65:30]
  assign cell_7_clock = clock;
  assign cell_7_reset = reset;
  assign cell_7_io_en = io_en; // @[act.scala 62:22]
  assign cell_7_io_i_data = io_i_data_7; // @[act.scala 63:26]
  assign cell_7_io_scale = io_scale; // @[act.scala 64:25]
  assign cell_7_io_zero_point = io_zero_point; // @[act.scala 65:30]
endmodule
module Calc_offset_0(
  input  [22:0] io_frac,
  output [4:0]  io_off
);
  wire [6:0] io_off_hi = io_frac[22:16]; // @[CircuitMath.scala 33:17]
  wire [15:0] io_off_lo = io_frac[15:0]; // @[CircuitMath.scala 34:17]
  wire  io_off_useHi = |io_off_hi; // @[CircuitMath.scala 35:22]
  wire [2:0] io_off_hi_1 = io_off_hi[6:4]; // @[CircuitMath.scala 33:17]
  wire [3:0] io_off_lo_1 = io_off_hi[3:0]; // @[CircuitMath.scala 34:17]
  wire  io_off_useHi_1 = |io_off_hi_1; // @[CircuitMath.scala 35:22]
  wire [1:0] _io_off_T_2 = io_off_hi_1[2] ? 2'h2 : {{1'd0}, io_off_hi_1[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_6 = io_off_lo_1[2] ? 2'h2 : {{1'd0}, io_off_lo_1[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_7 = io_off_lo_1[3] ? 2'h3 : _io_off_T_6; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_8 = io_off_useHi_1 ? _io_off_T_2 : _io_off_T_7; // @[CircuitMath.scala 36:21]
  wire [2:0] _io_off_T_9 = {io_off_useHi_1,_io_off_T_8}; // @[Cat.scala 33:92]
  wire [7:0] io_off_hi_2 = io_off_lo[15:8]; // @[CircuitMath.scala 33:17]
  wire [7:0] io_off_lo_2 = io_off_lo[7:0]; // @[CircuitMath.scala 34:17]
  wire  io_off_useHi_2 = |io_off_hi_2; // @[CircuitMath.scala 35:22]
  wire [3:0] io_off_hi_3 = io_off_hi_2[7:4]; // @[CircuitMath.scala 33:17]
  wire [3:0] io_off_lo_3 = io_off_hi_2[3:0]; // @[CircuitMath.scala 34:17]
  wire  io_off_useHi_3 = |io_off_hi_3; // @[CircuitMath.scala 35:22]
  wire [1:0] _io_off_T_13 = io_off_hi_3[2] ? 2'h2 : {{1'd0}, io_off_hi_3[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_14 = io_off_hi_3[3] ? 2'h3 : _io_off_T_13; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_18 = io_off_lo_3[2] ? 2'h2 : {{1'd0}, io_off_lo_3[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_19 = io_off_lo_3[3] ? 2'h3 : _io_off_T_18; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_20 = io_off_useHi_3 ? _io_off_T_14 : _io_off_T_19; // @[CircuitMath.scala 36:21]
  wire [2:0] _io_off_T_21 = {io_off_useHi_3,_io_off_T_20}; // @[Cat.scala 33:92]
  wire [3:0] io_off_hi_4 = io_off_lo_2[7:4]; // @[CircuitMath.scala 33:17]
  wire [3:0] io_off_lo_4 = io_off_lo_2[3:0]; // @[CircuitMath.scala 34:17]
  wire  io_off_useHi_4 = |io_off_hi_4; // @[CircuitMath.scala 35:22]
  wire [1:0] _io_off_T_25 = io_off_hi_4[2] ? 2'h2 : {{1'd0}, io_off_hi_4[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_26 = io_off_hi_4[3] ? 2'h3 : _io_off_T_25; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_30 = io_off_lo_4[2] ? 2'h2 : {{1'd0}, io_off_lo_4[1]}; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_31 = io_off_lo_4[3] ? 2'h3 : _io_off_T_30; // @[CircuitMath.scala 30:10]
  wire [1:0] _io_off_T_32 = io_off_useHi_4 ? _io_off_T_26 : _io_off_T_31; // @[CircuitMath.scala 36:21]
  wire [2:0] _io_off_T_33 = {io_off_useHi_4,_io_off_T_32}; // @[Cat.scala 33:92]
  wire [2:0] _io_off_T_34 = io_off_useHi_2 ? _io_off_T_21 : _io_off_T_33; // @[CircuitMath.scala 36:21]
  wire [3:0] _io_off_T_35 = {io_off_useHi_2,_io_off_T_34}; // @[Cat.scala 33:92]
  wire [3:0] _io_off_T_36 = io_off_useHi ? {{1'd0}, _io_off_T_9} : _io_off_T_35; // @[CircuitMath.scala 36:21]
  wire [4:0] _io_off_T_37 = {io_off_useHi,_io_off_T_36}; // @[Cat.scala 33:92]
  assign io_off = 5'h16 - _io_off_T_37; // @[FP32.scala 162:18]
endmodule
module FP32_Adder(
  input         clock,
  input         reset,
  input  [31:0] io_x,
  input  [31:0] io_y,
  output [31:0] io_z,
  input         io_valid_in
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [22:0] off0_io_frac; // @[FP32.scala 166:23]
  wire [4:0] off0_io_off; // @[FP32.scala 166:23]
  wire  xs_0 = io_x[31]; // @[FP32.scala 76:51]
  wire [7:0] xe_0 = io_x[30:23]; // @[FP32.scala 76:61]
  wire [22:0] xf_0 = io_x[22:0]; // @[FP32.scala 76:75]
  wire  ys_0 = io_y[31]; // @[FP32.scala 76:88]
  wire [7:0] ye_0 = io_y[30:23]; // @[FP32.scala 76:98]
  wire [22:0] yf_0 = io_y[22:0]; // @[FP32.scala 76:112]
  wire  y_gt_x_0 = io_y[30:0] > io_x[30:0]; // @[FP32.scala 79:30]
  wire [7:0] ze_0 = y_gt_x_0 ? ye_0 : xe_0; // @[FP32.scala 82:21]
  wire  _xf1_0_T = ye_0 != 8'h0; // @[FP32.scala 84:40]
  wire [23:0] _xf1_0_T_1 = {_xf1_0_T,yf_0}; // @[Cat.scala 33:92]
  wire  _xf1_0_T_2 = xe_0 != 8'h0; // @[FP32.scala 84:65]
  wire [23:0] _xf1_0_T_3 = {_xf1_0_T_2,xf_0}; // @[Cat.scala 33:92]
  wire [7:0] _xe_ye_0_T_1 = y_gt_x_0 ? xe_0 : ye_0; // @[FP32.scala 86:48]
  wire [7:0] xe_ye_0 = ze_0 - _xe_ye_0_T_1; // @[FP32.scala 86:43]
  reg  zs_a; // @[Reg.scala 19:16]
  reg [7:0] ze_a; // @[Reg.scala 19:16]
  reg [23:0] xf1_a; // @[Reg.scala 19:16]
  reg [23:0] yf1_a; // @[Reg.scala 19:16]
  reg [7:0] xe_ye_a; // @[Reg.scala 19:16]
  wire  _xs_ys_a_T = xs_0 == ys_0; // @[FP32.scala 93:32]
  reg  xs_ys_a; // @[Reg.scala 19:16]
  wire [4:0] xe_ye_reduced = xe_ye_a[4:0]; // @[FP32.scala 95:30]
  wire  xe_ye_32 = xe_ye_a[7:5] != 3'h0; // @[FP32.scala 96:37]
  wire [23:0] yf2_a0 = xe_ye_32 ? 24'h0 : yf1_a; // @[FP32.scala 97:26]
  wire [23:0] yf2_a1 = xe_ye_reduced[4] ? {{16'd0}, yf2_a0[23:16]} : yf2_a0; // @[FP32.scala 98:26]
  wire [23:0] yf2_a2 = xe_ye_reduced[3] ? {{8'd0}, yf2_a1[23:8]} : yf2_a1; // @[FP32.scala 99:26]
  wire [23:0] yf2_a3 = xe_ye_reduced[2] ? {{4'd0}, yf2_a2[23:4]} : yf2_a2; // @[FP32.scala 100:26]
  wire [23:0] yf2_a4 = xe_ye_reduced[1] ? {{2'd0}, yf2_a3[23:2]} : yf2_a3; // @[FP32.scala 101:26]
  reg  valid_1; // @[FP32.scala 104:24]
  reg  xs_ys_1; // @[Reg.scala 19:16]
  reg [23:0] xf1_1; // @[Reg.scala 19:16]
  reg [23:0] yf2_1; // @[Reg.scala 19:16]
  reg [7:0] ze_1; // @[Reg.scala 19:16]
  reg  zs_1; // @[Reg.scala 19:16]
  wire [24:0] _zf_1_T = xf1_1 + yf2_1; // @[FP32.scala 111:33]
  wire [23:0] _zf_1_T_2 = xf1_1 - yf2_1; // @[FP32.scala 111:49]
  reg  valid_2; // @[FP32.scala 113:24]
  reg [7:0] ze_2; // @[Reg.scala 19:16]
  reg  zs_2; // @[Reg.scala 19:16]
  reg [24:0] zf_2; // @[Reg.scala 19:16]
  reg  valid_3; // @[FP32.scala 122:25]
  reg [7:0] ze_3; // @[Reg.scala 19:16]
  reg  zs_3; // @[Reg.scala 19:16]
  reg [24:0] zf_3; // @[Reg.scala 19:16]
  reg [4:0] offset_3; // @[Reg.scala 19:16]
  wire [7:0] _GEN_19 = {{3'd0}, offset_3}; // @[FP32.scala 128:28]
  wire  underflow_3 = ze_3 < _GEN_19; // @[FP32.scala 128:28]
  wire  shift_right_3 = zf_3[24]; // @[FP32.scala 129:27]
  wire [7:0] _ze1_3_T_1 = ze_3 + 8'h1; // @[FP32.scala 133:30]
  wire [7:0] _ze1_3_T_3 = ze_3 - _GEN_19; // @[FP32.scala 134:23]
  wire [7:0] _ze1_3_T_4 = shift_right_3 ? _ze1_3_T_1 : _ze1_3_T_3; // @[Mux.scala 47:70]
  wire [7:0] ze1_3 = underflow_3 ? 8'h0 : _ze1_3_T_4; // @[Mux.scala 47:70]
  wire [55:0] _GEN_0 = {{31'd0}, zf_3}; // @[FP32.scala 141:23]
  wire [55:0] _zf1_3_T_1 = _GEN_0 << offset_3; // @[FP32.scala 141:23]
  wire [22:0] _zf1_3_T_3 = shift_right_3 ? zf_3[23:1] : _zf1_3_T_1[22:0]; // @[Mux.scala 47:70]
  wire [22:0] zf1_3 = underflow_3 ? 23'h0 : _zf1_3_T_3; // @[Mux.scala 47:70]
  reg  valid_4; // @[FP32.scala 146:24]
  wire [31:0] _io_z_T = {zs_3,ze1_3,zf1_3}; // @[Cat.scala 33:92]
  reg [31:0] io_z_r; // @[Reg.scala 19:16]
  Calc_offset_0 off0 ( // @[FP32.scala 166:23]
    .io_frac(off0_io_frac),
    .io_off(off0_io_off)
  );
  assign io_z = io_z_r; // @[FP32.scala 147:8]
  assign off0_io_frac = zf_2[23:1]; // @[FP32.scala 118:23]
  always @(posedge clock) begin
    if (io_valid_in) begin // @[Reg.scala 20:18]
      if (y_gt_x_0) begin // @[FP32.scala 81:21]
        zs_a <= ys_0;
      end else begin
        zs_a <= xs_0;
      end
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      if (y_gt_x_0) begin // @[FP32.scala 82:21]
        ze_a <= ye_0;
      end else begin
        ze_a <= xe_0;
      end
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      if (y_gt_x_0) begin // @[FP32.scala 84:20]
        xf1_a <= _xf1_0_T_1;
      end else begin
        xf1_a <= _xf1_0_T_3;
      end
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      if (y_gt_x_0) begin // @[FP32.scala 85:20]
        yf1_a <= _xf1_0_T_3;
      end else begin
        yf1_a <= _xf1_0_T_1;
      end
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      xe_ye_a <= xe_ye_0; // @[Reg.scala 20:22]
    end
    if (io_valid_in) begin // @[Reg.scala 20:18]
      xs_ys_a <= _xs_ys_a_T; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[FP32.scala 104:24]
      valid_1 <= 1'h0; // @[FP32.scala 104:24]
    end else begin
      valid_1 <= io_valid_in; // @[FP32.scala 104:24]
    end
    if (valid_1) begin // @[Reg.scala 20:18]
      xs_ys_1 <= xs_ys_a; // @[Reg.scala 20:22]
    end
    if (valid_1) begin // @[Reg.scala 20:18]
      xf1_1 <= xf1_a; // @[Reg.scala 20:22]
    end
    if (valid_1) begin // @[Reg.scala 20:18]
      if (xe_ye_reduced[0]) begin // @[FP32.scala 102:26]
        yf2_1 <= {{1'd0}, yf2_a4[23:1]};
      end else if (xe_ye_reduced[1]) begin // @[FP32.scala 101:26]
        yf2_1 <= {{2'd0}, yf2_a3[23:2]};
      end else if (xe_ye_reduced[2]) begin // @[FP32.scala 100:26]
        yf2_1 <= {{4'd0}, yf2_a2[23:4]};
      end else begin
        yf2_1 <= yf2_a2;
      end
    end
    if (valid_1) begin // @[Reg.scala 20:18]
      ze_1 <= ze_a; // @[Reg.scala 20:22]
    end
    if (valid_1) begin // @[Reg.scala 20:18]
      zs_1 <= zs_a; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[FP32.scala 113:24]
      valid_2 <= 1'h0; // @[FP32.scala 113:24]
    end else begin
      valid_2 <= valid_1; // @[FP32.scala 113:24]
    end
    if (valid_2) begin // @[Reg.scala 20:18]
      ze_2 <= ze_1; // @[Reg.scala 20:22]
    end
    if (valid_2) begin // @[Reg.scala 20:18]
      zs_2 <= zs_1; // @[Reg.scala 20:22]
    end
    if (valid_2) begin // @[Reg.scala 20:18]
      if (xs_ys_1) begin // @[FP32.scala 111:17]
        zf_2 <= _zf_1_T;
      end else begin
        zf_2 <= {{1'd0}, _zf_1_T_2};
      end
    end
    if (reset) begin // @[FP32.scala 122:25]
      valid_3 <= 1'h0; // @[FP32.scala 122:25]
    end else begin
      valid_3 <= valid_2; // @[FP32.scala 122:25]
    end
    if (valid_3) begin // @[Reg.scala 20:18]
      ze_3 <= ze_2; // @[Reg.scala 20:22]
    end
    if (valid_3) begin // @[Reg.scala 20:18]
      zs_3 <= zs_2; // @[Reg.scala 20:22]
    end
    if (valid_3) begin // @[Reg.scala 20:18]
      zf_3 <= zf_2; // @[Reg.scala 20:22]
    end
    if (valid_3) begin // @[Reg.scala 20:18]
      offset_3 <= off0_io_off; // @[Reg.scala 20:22]
    end
    if (reset) begin // @[FP32.scala 146:24]
      valid_4 <= 1'h0; // @[FP32.scala 146:24]
    end else begin
      valid_4 <= valid_3; // @[FP32.scala 146:24]
    end
    if (valid_4) begin // @[Reg.scala 20:18]
      io_z_r <= _io_z_T; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  zs_a = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ze_a = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  xf1_a = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  yf1_a = _RAND_3[23:0];
  _RAND_4 = {1{`RANDOM}};
  xe_ye_a = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  xs_ys_a = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  valid_1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  xs_ys_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  xf1_1 = _RAND_8[23:0];
  _RAND_9 = {1{`RANDOM}};
  yf2_1 = _RAND_9[23:0];
  _RAND_10 = {1{`RANDOM}};
  ze_1 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  zs_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  valid_2 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  ze_2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  zs_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  zf_2 = _RAND_15[24:0];
  _RAND_16 = {1{`RANDOM}};
  valid_3 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ze_3 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  zs_3 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  zf_3 = _RAND_19[24:0];
  _RAND_20 = {1{`RANDOM}};
  offset_3 = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  valid_4 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  io_z_r = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cal_add_zero_point(
  input        clock,
  input        reset,
  input  [7:0] io_zero_point,
  input  [7:0] io_data_in,
  output [7:0] io_data_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] out; // @[quant.scala 107:22]
  wire [7:0] _out_T_2 = $signed(io_data_in) + $signed(io_zero_point); // @[quant.scala 108:15]
  assign io_data_out = out; // @[quant.scala 109:24]
  always @(posedge clock) begin
    if (reset) begin // @[quant.scala 107:22]
      out <= 8'sh0; // @[quant.scala 107:22]
    end else begin
      out <= _out_T_2; // @[quant.scala 108:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RecFNToIN_e8_s24_i8(
  input  [32:0] io_in,
  output [7:0]  io_out
);
  wire [8:0] rawIn_exp = io_in[31:23]; // @[rawFloatFromRecFN.scala 50:21]
  wire  rawIn_isZero = rawIn_exp[8:6] == 3'h0; // @[rawFloatFromRecFN.scala 51:53]
  wire  rawIn_isSpecial = rawIn_exp[8:7] == 2'h3; // @[rawFloatFromRecFN.scala 52:53]
  wire  rawIn__isNaN = rawIn_isSpecial & rawIn_exp[6]; // @[rawFloatFromRecFN.scala 55:33]
  wire  rawIn__isInf = rawIn_isSpecial & ~rawIn_exp[6]; // @[rawFloatFromRecFN.scala 56:33]
  wire  rawIn__sign = io_in[32]; // @[rawFloatFromRecFN.scala 58:25]
  wire [9:0] rawIn__sExp = {1'b0,$signed(rawIn_exp)}; // @[rawFloatFromRecFN.scala 59:27]
  wire  _rawIn_out_sig_T = ~rawIn_isZero; // @[rawFloatFromRecFN.scala 60:35]
  wire [24:0] rawIn__sig = {1'h0,_rawIn_out_sig_T,io_in[22:0]}; // @[rawFloatFromRecFN.scala 60:44]
  wire  magGeOne = rawIn__sExp[8]; // @[RecFNToIN.scala 61:30]
  wire [7:0] posExp = rawIn__sExp[7:0]; // @[RecFNToIN.scala 62:28]
  wire  magJustBelowOne = ~magGeOne & &posExp; // @[RecFNToIN.scala 63:37]
  wire [23:0] _shiftedSig_T_1 = {magGeOne,rawIn__sig[22:0]}; // @[RecFNToIN.scala 83:19]
  wire [2:0] _shiftedSig_T_3 = magGeOne ? rawIn__sExp[2:0] : 3'h0; // @[RecFNToIN.scala 84:16]
  wire [30:0] _GEN_1 = {{7'd0}, _shiftedSig_T_1}; // @[RecFNToIN.scala 83:49]
  wire [30:0] shiftedSig = _GEN_1 << _shiftedSig_T_3; // @[RecFNToIN.scala 83:49]
  wire [9:0] alignedSig = {shiftedSig[30:22],|shiftedSig[21:0]}; // @[RecFNToIN.scala 89:38]
  wire [7:0] unroundedInt = alignedSig[9:2]; // @[RecFNToIN.scala 90:52]
  wire  roundIncr_near_maxMag = magGeOne & alignedSig[1] | magJustBelowOne; // @[RecFNToIN.scala 96:61]
  wire [7:0] _complUnroundedInt_T = ~unroundedInt; // @[RecFNToIN.scala 103:45]
  wire [7:0] complUnroundedInt = rawIn__sign ? _complUnroundedInt_T : unroundedInt; // @[RecFNToIN.scala 103:32]
  wire [7:0] _roundedInt_T_2 = complUnroundedInt + 8'h1; // @[RecFNToIN.scala 106:31]
  wire [7:0] roundedInt = roundIncr_near_maxMag ^ rawIn__sign ? _roundedInt_T_2 : complUnroundedInt; // @[RecFNToIN.scala 105:12]
  wire  magGeOne_atOverflowEdge = posExp == 8'h7; // @[RecFNToIN.scala 110:43]
  wire  roundCarryBut2 = &unroundedInt[5:0] & roundIncr_near_maxMag; // @[RecFNToIN.scala 113:61]
  wire  _common_overflow_T_3 = |unroundedInt[6:0] | roundIncr_near_maxMag; // @[RecFNToIN.scala 120:64]
  wire  _common_overflow_T_4 = magGeOne_atOverflowEdge & _common_overflow_T_3; // @[RecFNToIN.scala 119:49]
  wire  _common_overflow_T_6 = posExp == 8'h6 & roundCarryBut2; // @[RecFNToIN.scala 122:60]
  wire  _common_overflow_T_7 = magGeOne_atOverflowEdge | _common_overflow_T_6; // @[RecFNToIN.scala 121:49]
  wire  _common_overflow_T_8 = rawIn__sign ? _common_overflow_T_4 : _common_overflow_T_7; // @[RecFNToIN.scala 118:24]
  wire  _common_overflow_T_14 = posExp >= 8'h8 | _common_overflow_T_8; // @[RecFNToIN.scala 116:36]
  wire  common_overflow = magGeOne & _common_overflow_T_14; // @[RecFNToIN.scala 115:12]
  wire  invalidExc = rawIn__isNaN | rawIn__isInf; // @[RecFNToIN.scala 133:34]
  wire  excSign = ~rawIn__isNaN & rawIn__sign; // @[RecFNToIN.scala 137:32]
  wire [7:0] _excOut_T_1 = excSign ? 8'h80 : 8'h0; // @[RecFNToIN.scala 139:12]
  wire [6:0] _excOut_T_3 = ~excSign ? 7'h7f : 7'h0; // @[RecFNToIN.scala 143:12]
  wire [7:0] _GEN_0 = {{1'd0}, _excOut_T_3}; // @[RecFNToIN.scala 142:11]
  wire [7:0] excOut = _excOut_T_1 | _GEN_0; // @[RecFNToIN.scala 142:11]
  assign io_out = invalidExc | common_overflow ? excOut : roundedInt; // @[RecFNToIN.scala 145:18]
endmodule
module quant_cell(
  input         clock,
  input         reset,
  input         io_en,
  input  [31:0] io_i_data,
  input  [31:0] io_scale,
  output [7:0]  io_o_data,
  input  [7:0]  io_zero_point
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  add_module_clock; // @[act.scala 203:28]
  wire  add_module_reset; // @[act.scala 203:28]
  wire [7:0] add_module_io_zero_point; // @[act.scala 203:28]
  wire [7:0] add_module_io_data_in; // @[act.scala 203:28]
  wire [7:0] add_module_io_data_out; // @[act.scala 203:28]
  wire  quant_data_muler_clock; // @[Arithmetic.scala 95:25]
  wire  quant_data_muler_reset; // @[Arithmetic.scala 95:25]
  wire [31:0] quant_data_muler_io_x; // @[Arithmetic.scala 95:25]
  wire [31:0] quant_data_muler_io_y; // @[Arithmetic.scala 95:25]
  wire [31:0] quant_data_muler_io_z; // @[Arithmetic.scala 95:25]
  wire  quant_data_muler_io_valid_in; // @[Arithmetic.scala 95:25]
  wire [32:0] add_in_convert_io_in; // @[Arithmetic.scala 60:25]
  wire [7:0] add_in_convert_io_out; // @[Arithmetic.scala 60:25]
  reg [31:0] i_data_t; // @[Reg.scala 35:20]
  wire [31:0] quant_data_bits = quant_data_muler_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire  add_in_convert_io_in_rawIn_sign = quant_data_bits[31]; // @[rawFloatFromFN.scala 44:18]
  wire [7:0] add_in_convert_io_in_rawIn_expIn = quant_data_bits[30:23]; // @[rawFloatFromFN.scala 45:19]
  wire [22:0] add_in_convert_io_in_rawIn_fractIn = quant_data_bits[22:0]; // @[rawFloatFromFN.scala 46:21]
  wire  add_in_convert_io_in_rawIn_isZeroExpIn = add_in_convert_io_in_rawIn_expIn == 8'h0; // @[rawFloatFromFN.scala 48:30]
  wire  add_in_convert_io_in_rawIn_isZeroFractIn = add_in_convert_io_in_rawIn_fractIn == 23'h0; // @[rawFloatFromFN.scala 49:34]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_23 = add_in_convert_io_in_rawIn_fractIn[1] ? 5'h15 : 5'h16; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_24 = add_in_convert_io_in_rawIn_fractIn[2] ? 5'h14 :
    _add_in_convert_io_in_rawIn_normDist_T_23; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_25 = add_in_convert_io_in_rawIn_fractIn[3] ? 5'h13 :
    _add_in_convert_io_in_rawIn_normDist_T_24; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_26 = add_in_convert_io_in_rawIn_fractIn[4] ? 5'h12 :
    _add_in_convert_io_in_rawIn_normDist_T_25; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_27 = add_in_convert_io_in_rawIn_fractIn[5] ? 5'h11 :
    _add_in_convert_io_in_rawIn_normDist_T_26; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_28 = add_in_convert_io_in_rawIn_fractIn[6] ? 5'h10 :
    _add_in_convert_io_in_rawIn_normDist_T_27; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_29 = add_in_convert_io_in_rawIn_fractIn[7] ? 5'hf :
    _add_in_convert_io_in_rawIn_normDist_T_28; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_30 = add_in_convert_io_in_rawIn_fractIn[8] ? 5'he :
    _add_in_convert_io_in_rawIn_normDist_T_29; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_31 = add_in_convert_io_in_rawIn_fractIn[9] ? 5'hd :
    _add_in_convert_io_in_rawIn_normDist_T_30; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_32 = add_in_convert_io_in_rawIn_fractIn[10] ? 5'hc :
    _add_in_convert_io_in_rawIn_normDist_T_31; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_33 = add_in_convert_io_in_rawIn_fractIn[11] ? 5'hb :
    _add_in_convert_io_in_rawIn_normDist_T_32; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_34 = add_in_convert_io_in_rawIn_fractIn[12] ? 5'ha :
    _add_in_convert_io_in_rawIn_normDist_T_33; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_35 = add_in_convert_io_in_rawIn_fractIn[13] ? 5'h9 :
    _add_in_convert_io_in_rawIn_normDist_T_34; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_36 = add_in_convert_io_in_rawIn_fractIn[14] ? 5'h8 :
    _add_in_convert_io_in_rawIn_normDist_T_35; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_37 = add_in_convert_io_in_rawIn_fractIn[15] ? 5'h7 :
    _add_in_convert_io_in_rawIn_normDist_T_36; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_38 = add_in_convert_io_in_rawIn_fractIn[16] ? 5'h6 :
    _add_in_convert_io_in_rawIn_normDist_T_37; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_39 = add_in_convert_io_in_rawIn_fractIn[17] ? 5'h5 :
    _add_in_convert_io_in_rawIn_normDist_T_38; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_40 = add_in_convert_io_in_rawIn_fractIn[18] ? 5'h4 :
    _add_in_convert_io_in_rawIn_normDist_T_39; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_41 = add_in_convert_io_in_rawIn_fractIn[19] ? 5'h3 :
    _add_in_convert_io_in_rawIn_normDist_T_40; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_42 = add_in_convert_io_in_rawIn_fractIn[20] ? 5'h2 :
    _add_in_convert_io_in_rawIn_normDist_T_41; // @[Mux.scala 47:70]
  wire [4:0] _add_in_convert_io_in_rawIn_normDist_T_43 = add_in_convert_io_in_rawIn_fractIn[21] ? 5'h1 :
    _add_in_convert_io_in_rawIn_normDist_T_42; // @[Mux.scala 47:70]
  wire [4:0] add_in_convert_io_in_rawIn_normDist = add_in_convert_io_in_rawIn_fractIn[22] ? 5'h0 :
    _add_in_convert_io_in_rawIn_normDist_T_43; // @[Mux.scala 47:70]
  wire [53:0] _GEN_2 = {{31'd0}, add_in_convert_io_in_rawIn_fractIn}; // @[rawFloatFromFN.scala 52:33]
  wire [53:0] _add_in_convert_io_in_rawIn_subnormFract_T = _GEN_2 << add_in_convert_io_in_rawIn_normDist; // @[rawFloatFromFN.scala 52:33]
  wire [22:0] add_in_convert_io_in_rawIn_subnormFract = {_add_in_convert_io_in_rawIn_subnormFract_T[21:0], 1'h0}; // @[rawFloatFromFN.scala 52:64]
  wire [8:0] _GEN_3 = {{4'd0}, add_in_convert_io_in_rawIn_normDist}; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _add_in_convert_io_in_rawIn_adjustedExp_T = _GEN_3 ^ 9'h1ff; // @[rawFloatFromFN.scala 55:18]
  wire [8:0] _add_in_convert_io_in_rawIn_adjustedExp_T_1 = add_in_convert_io_in_rawIn_isZeroExpIn ?
    _add_in_convert_io_in_rawIn_adjustedExp_T : {{1'd0}, add_in_convert_io_in_rawIn_expIn}; // @[rawFloatFromFN.scala 54:10]
  wire [1:0] _add_in_convert_io_in_rawIn_adjustedExp_T_2 = add_in_convert_io_in_rawIn_isZeroExpIn ? 2'h2 : 2'h1; // @[rawFloatFromFN.scala 58:14]
  wire [7:0] _GEN_4 = {{6'd0}, _add_in_convert_io_in_rawIn_adjustedExp_T_2}; // @[rawFloatFromFN.scala 58:9]
  wire [7:0] _add_in_convert_io_in_rawIn_adjustedExp_T_3 = 8'h80 | _GEN_4; // @[rawFloatFromFN.scala 58:9]
  wire [8:0] _GEN_5 = {{1'd0}, _add_in_convert_io_in_rawIn_adjustedExp_T_3}; // @[rawFloatFromFN.scala 57:9]
  wire [8:0] add_in_convert_io_in_rawIn_adjustedExp = _add_in_convert_io_in_rawIn_adjustedExp_T_1 + _GEN_5; // @[rawFloatFromFN.scala 57:9]
  wire  add_in_convert_io_in_rawIn_isZero = add_in_convert_io_in_rawIn_isZeroExpIn &
    add_in_convert_io_in_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 60:30]
  wire  add_in_convert_io_in_rawIn_isSpecial = add_in_convert_io_in_rawIn_adjustedExp[8:7] == 2'h3; // @[rawFloatFromFN.scala 61:57]
  wire  add_in_convert_io_in_rawIn__isNaN = add_in_convert_io_in_rawIn_isSpecial & ~
    add_in_convert_io_in_rawIn_isZeroFractIn; // @[rawFloatFromFN.scala 64:28]
  wire [9:0] add_in_convert_io_in_rawIn__sExp = {1'b0,$signed(add_in_convert_io_in_rawIn_adjustedExp)}; // @[rawFloatFromFN.scala 68:42]
  wire  _add_in_convert_io_in_rawIn_out_sig_T = ~add_in_convert_io_in_rawIn_isZero; // @[rawFloatFromFN.scala 70:19]
  wire [22:0] _add_in_convert_io_in_rawIn_out_sig_T_2 = add_in_convert_io_in_rawIn_isZeroExpIn ?
    add_in_convert_io_in_rawIn_subnormFract : add_in_convert_io_in_rawIn_fractIn; // @[rawFloatFromFN.scala 70:33]
  wire [24:0] add_in_convert_io_in_rawIn__sig = {1'h0,_add_in_convert_io_in_rawIn_out_sig_T,
    _add_in_convert_io_in_rawIn_out_sig_T_2}; // @[rawFloatFromFN.scala 70:27]
  wire [2:0] _add_in_convert_io_in_T_1 = add_in_convert_io_in_rawIn_isZero ? 3'h0 : add_in_convert_io_in_rawIn__sExp[8:6
    ]; // @[recFNFromFN.scala 48:15]
  wire [2:0] _GEN_6 = {{2'd0}, add_in_convert_io_in_rawIn__isNaN}; // @[recFNFromFN.scala 48:76]
  wire [2:0] _add_in_convert_io_in_T_3 = _add_in_convert_io_in_T_1 | _GEN_6; // @[recFNFromFN.scala 48:76]
  wire [9:0] _add_in_convert_io_in_T_6 = {add_in_convert_io_in_rawIn_sign,_add_in_convert_io_in_T_3,
    add_in_convert_io_in_rawIn__sExp[5:0]}; // @[recFNFromFN.scala 49:45]
  reg [7:0] add_in_res; // @[Reg.scala 35:20]
  reg  add_in_REG; // @[Arithmetic.scala 65:66]
  reg [7:0] add_in_r; // @[Reg.scala 19:16]
  cal_add_zero_point add_module ( // @[act.scala 203:28]
    .clock(add_module_clock),
    .reset(add_module_reset),
    .io_zero_point(add_module_io_zero_point),
    .io_data_in(add_module_io_data_in),
    .io_data_out(add_module_io_data_out)
  );
  FP32_Mult quant_data_muler ( // @[Arithmetic.scala 95:25]
    .clock(quant_data_muler_clock),
    .reset(quant_data_muler_reset),
    .io_x(quant_data_muler_io_x),
    .io_y(quant_data_muler_io_y),
    .io_z(quant_data_muler_io_z),
    .io_valid_in(quant_data_muler_io_valid_in)
  );
  RecFNToIN_e8_s24_i8 add_in_convert ( // @[Arithmetic.scala 60:25]
    .io_in(add_in_convert_io_in),
    .io_out(add_in_convert_io_out)
  );
  assign io_o_data = add_module_io_data_out; // @[act.scala 206:15]
  assign add_module_clock = clock;
  assign add_module_reset = reset;
  assign add_module_io_zero_point = io_zero_point; // @[act.scala 204:30]
  assign add_module_io_data_in = add_in_r; // @[act.scala 209:55]
  assign quant_data_muler_clock = clock;
  assign quant_data_muler_reset = reset;
  assign quant_data_muler_io_x = i_data_t; // @[Arithmetic.scala 124:22 125:17]
  assign quant_data_muler_io_y = io_scale; // @[Arithmetic.scala 124:22 125:17]
  assign quant_data_muler_io_valid_in = io_en; // @[Arithmetic.scala 98:25]
  assign add_in_convert_io_in = {_add_in_convert_io_in_T_6,add_in_convert_io_in_rawIn__sig[22:0]}; // @[recFNFromFN.scala 50:41]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      i_data_t <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      i_data_t <= io_i_data; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      add_in_res <= 8'sh0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      add_in_res <= add_in_convert_io_out; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Arithmetic.scala 65:66]
      add_in_REG <= 1'h0; // @[Arithmetic.scala 65:66]
    end else begin
      add_in_REG <= io_en; // @[Arithmetic.scala 65:66]
    end
    if (add_in_REG) begin // @[Reg.scala 20:18]
      if ($signed(add_in_res) == 8'sh80) begin // @[Arithmetic.scala 65:18]
        add_in_r <= -8'sh7f;
      end else begin
        add_in_r <= add_in_res;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_data_t = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  add_in_res = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  add_in_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  add_in_r = _RAND_3[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module quant_fp32_2_int8(
  input         clock,
  input         reset,
  input         io_en,
  input  [31:0] io_i_data_0,
  input  [31:0] io_i_data_1,
  input  [31:0] io_i_data_2,
  input  [31:0] io_i_data_3,
  input  [31:0] io_i_data_4,
  input  [31:0] io_i_data_5,
  input  [31:0] io_i_data_6,
  input  [31:0] io_i_data_7,
  input  [31:0] io_scale,
  input  [7:0]  io_zero_point,
  output [7:0]  io_o_data_0,
  output [7:0]  io_o_data_1,
  output [7:0]  io_o_data_2,
  output [7:0]  io_o_data_3,
  output [7:0]  io_o_data_4,
  output [7:0]  io_o_data_5,
  output [7:0]  io_o_data_6,
  output [7:0]  io_o_data_7
);
  wire  cell_0_clock; // @[act.scala 38:36]
  wire  cell_0_reset; // @[act.scala 38:36]
  wire  cell_0_io_en; // @[act.scala 38:36]
  wire [31:0] cell_0_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_0_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_0_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_0_io_zero_point; // @[act.scala 38:36]
  wire  cell_1_clock; // @[act.scala 38:36]
  wire  cell_1_reset; // @[act.scala 38:36]
  wire  cell_1_io_en; // @[act.scala 38:36]
  wire [31:0] cell_1_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_1_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_1_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_1_io_zero_point; // @[act.scala 38:36]
  wire  cell_2_clock; // @[act.scala 38:36]
  wire  cell_2_reset; // @[act.scala 38:36]
  wire  cell_2_io_en; // @[act.scala 38:36]
  wire [31:0] cell_2_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_2_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_2_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_2_io_zero_point; // @[act.scala 38:36]
  wire  cell_3_clock; // @[act.scala 38:36]
  wire  cell_3_reset; // @[act.scala 38:36]
  wire  cell_3_io_en; // @[act.scala 38:36]
  wire [31:0] cell_3_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_3_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_3_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_3_io_zero_point; // @[act.scala 38:36]
  wire  cell_4_clock; // @[act.scala 38:36]
  wire  cell_4_reset; // @[act.scala 38:36]
  wire  cell_4_io_en; // @[act.scala 38:36]
  wire [31:0] cell_4_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_4_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_4_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_4_io_zero_point; // @[act.scala 38:36]
  wire  cell_5_clock; // @[act.scala 38:36]
  wire  cell_5_reset; // @[act.scala 38:36]
  wire  cell_5_io_en; // @[act.scala 38:36]
  wire [31:0] cell_5_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_5_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_5_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_5_io_zero_point; // @[act.scala 38:36]
  wire  cell_6_clock; // @[act.scala 38:36]
  wire  cell_6_reset; // @[act.scala 38:36]
  wire  cell_6_io_en; // @[act.scala 38:36]
  wire [31:0] cell_6_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_6_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_6_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_6_io_zero_point; // @[act.scala 38:36]
  wire  cell_7_clock; // @[act.scala 38:36]
  wire  cell_7_reset; // @[act.scala 38:36]
  wire  cell_7_io_en; // @[act.scala 38:36]
  wire [31:0] cell_7_io_i_data; // @[act.scala 38:36]
  wire [31:0] cell_7_io_scale; // @[act.scala 38:36]
  wire [7:0] cell_7_io_o_data; // @[act.scala 38:36]
  wire [7:0] cell_7_io_zero_point; // @[act.scala 38:36]
  quant_cell cell_0 ( // @[act.scala 38:36]
    .clock(cell_0_clock),
    .reset(cell_0_reset),
    .io_en(cell_0_io_en),
    .io_i_data(cell_0_io_i_data),
    .io_scale(cell_0_io_scale),
    .io_o_data(cell_0_io_o_data),
    .io_zero_point(cell_0_io_zero_point)
  );
  quant_cell cell_1 ( // @[act.scala 38:36]
    .clock(cell_1_clock),
    .reset(cell_1_reset),
    .io_en(cell_1_io_en),
    .io_i_data(cell_1_io_i_data),
    .io_scale(cell_1_io_scale),
    .io_o_data(cell_1_io_o_data),
    .io_zero_point(cell_1_io_zero_point)
  );
  quant_cell cell_2 ( // @[act.scala 38:36]
    .clock(cell_2_clock),
    .reset(cell_2_reset),
    .io_en(cell_2_io_en),
    .io_i_data(cell_2_io_i_data),
    .io_scale(cell_2_io_scale),
    .io_o_data(cell_2_io_o_data),
    .io_zero_point(cell_2_io_zero_point)
  );
  quant_cell cell_3 ( // @[act.scala 38:36]
    .clock(cell_3_clock),
    .reset(cell_3_reset),
    .io_en(cell_3_io_en),
    .io_i_data(cell_3_io_i_data),
    .io_scale(cell_3_io_scale),
    .io_o_data(cell_3_io_o_data),
    .io_zero_point(cell_3_io_zero_point)
  );
  quant_cell cell_4 ( // @[act.scala 38:36]
    .clock(cell_4_clock),
    .reset(cell_4_reset),
    .io_en(cell_4_io_en),
    .io_i_data(cell_4_io_i_data),
    .io_scale(cell_4_io_scale),
    .io_o_data(cell_4_io_o_data),
    .io_zero_point(cell_4_io_zero_point)
  );
  quant_cell cell_5 ( // @[act.scala 38:36]
    .clock(cell_5_clock),
    .reset(cell_5_reset),
    .io_en(cell_5_io_en),
    .io_i_data(cell_5_io_i_data),
    .io_scale(cell_5_io_scale),
    .io_o_data(cell_5_io_o_data),
    .io_zero_point(cell_5_io_zero_point)
  );
  quant_cell cell_6 ( // @[act.scala 38:36]
    .clock(cell_6_clock),
    .reset(cell_6_reset),
    .io_en(cell_6_io_en),
    .io_i_data(cell_6_io_i_data),
    .io_scale(cell_6_io_scale),
    .io_o_data(cell_6_io_o_data),
    .io_zero_point(cell_6_io_zero_point)
  );
  quant_cell cell_7 ( // @[act.scala 38:36]
    .clock(cell_7_clock),
    .reset(cell_7_reset),
    .io_en(cell_7_io_en),
    .io_i_data(cell_7_io_i_data),
    .io_scale(cell_7_io_scale),
    .io_o_data(cell_7_io_o_data),
    .io_zero_point(cell_7_io_zero_point)
  );
  assign io_o_data_0 = cell_0_io_o_data; // @[act.scala 44:21]
  assign io_o_data_1 = cell_1_io_o_data; // @[act.scala 44:21]
  assign io_o_data_2 = cell_2_io_o_data; // @[act.scala 44:21]
  assign io_o_data_3 = cell_3_io_o_data; // @[act.scala 44:21]
  assign io_o_data_4 = cell_4_io_o_data; // @[act.scala 44:21]
  assign io_o_data_5 = cell_5_io_o_data; // @[act.scala 44:21]
  assign io_o_data_6 = cell_6_io_o_data; // @[act.scala 44:21]
  assign io_o_data_7 = cell_7_io_o_data; // @[act.scala 44:21]
  assign cell_0_clock = clock;
  assign cell_0_reset = reset;
  assign cell_0_io_en = io_en; // @[act.scala 40:22]
  assign cell_0_io_i_data = io_i_data_0; // @[act.scala 41:26]
  assign cell_0_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_0_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_1_clock = clock;
  assign cell_1_reset = reset;
  assign cell_1_io_en = io_en; // @[act.scala 40:22]
  assign cell_1_io_i_data = io_i_data_1; // @[act.scala 41:26]
  assign cell_1_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_1_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_2_clock = clock;
  assign cell_2_reset = reset;
  assign cell_2_io_en = io_en; // @[act.scala 40:22]
  assign cell_2_io_i_data = io_i_data_2; // @[act.scala 41:26]
  assign cell_2_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_2_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_3_clock = clock;
  assign cell_3_reset = reset;
  assign cell_3_io_en = io_en; // @[act.scala 40:22]
  assign cell_3_io_i_data = io_i_data_3; // @[act.scala 41:26]
  assign cell_3_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_3_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_4_clock = clock;
  assign cell_4_reset = reset;
  assign cell_4_io_en = io_en; // @[act.scala 40:22]
  assign cell_4_io_i_data = io_i_data_4; // @[act.scala 41:26]
  assign cell_4_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_4_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_5_clock = clock;
  assign cell_5_reset = reset;
  assign cell_5_io_en = io_en; // @[act.scala 40:22]
  assign cell_5_io_i_data = io_i_data_5; // @[act.scala 41:26]
  assign cell_5_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_5_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_6_clock = clock;
  assign cell_6_reset = reset;
  assign cell_6_io_en = io_en; // @[act.scala 40:22]
  assign cell_6_io_i_data = io_i_data_6; // @[act.scala 41:26]
  assign cell_6_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_6_io_zero_point = io_zero_point; // @[act.scala 43:30]
  assign cell_7_clock = clock;
  assign cell_7_reset = reset;
  assign cell_7_io_en = io_en; // @[act.scala 40:22]
  assign cell_7_io_i_data = io_i_data_7; // @[act.scala 41:26]
  assign cell_7_io_scale = io_scale; // @[act.scala 42:25]
  assign cell_7_io_zero_point = io_zero_point; // @[act.scala 43:30]
endmodule
module alu_act_param_select(
  input  [1:0]  io_act_op,
  output [31:0] io_cfg_act_coefficient_a_0,
  output [31:0] io_cfg_act_coefficient_a_1,
  output [31:0] io_cfg_act_coefficient_a_2,
  output [31:0] io_cfg_act_coefficient_a_3,
  output [31:0] io_cfg_act_coefficient_b_0,
  output [31:0] io_cfg_act_coefficient_b_1,
  output [31:0] io_cfg_act_coefficient_b_2,
  output [31:0] io_cfg_act_coefficient_b_3,
  output [31:0] io_cfg_act_coefficient_b_4,
  output [31:0] io_cfg_act_coefficient_c_0,
  output [31:0] io_cfg_act_coefficient_c_1,
  output [31:0] io_cfg_act_coefficient_c_2,
  output [31:0] io_cfg_act_coefficient_c_3,
  output [31:0] io_cfg_act_coefficient_c_4,
  output [31:0] io_cfg_act_range_0,
  output [31:0] io_cfg_act_range_1,
  output [31:0] io_cfg_act_range_2,
  output [31:0] io_cfg_act_range_3,
  output [1:0]  io_cfg_act_func_prop
);
  wire  act_op_sel_0 = io_act_op == 2'h0; // @[act.scala 173:70]
  wire  act_op_sel_1 = io_act_op == 2'h1; // @[act.scala 173:70]
  wire  act_op_sel_2 = io_act_op == 2'h2; // @[act.scala 173:70]
  wire [31:0] _act_coefficient_a_0_T = act_op_sel_2 ? 32'hbce448c5 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_0_T_1 = act_op_sel_1 ? 32'h0 : _act_coefficient_a_0_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_0_T = act_op_sel_2 ? 32'h3e855f24 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_0_T_1 = act_op_sel_1 ? 32'h0 : _act_coefficient_b_0_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_0_T = act_op_sel_2 ? 32'h3eff9198 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_0_T_1 = act_op_sel_1 ? 32'h0 : _act_coefficient_c_0_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_1_T = act_op_sel_2 ? 32'hbd3f460c : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_1_T_1 = act_op_sel_1 ? 32'hbc23b9f9 : _act_coefficient_a_1_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_1_T = act_op_sel_2 ? 32'h3e94471d : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_1_T_1 = act_op_sel_1 ? 32'hbe0aaa59 : _act_coefficient_b_1_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_1_T = act_op_sel_2 ? 32'h3ef9f7f8 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_1_T_1 = act_op_sel_1 ? 32'hbeebfcc8 : _act_coefficient_c_1_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_2_T = act_op_sel_2 ? 32'hbc718b08 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_2_T_1 = act_op_sel_1 ? 32'h3e490809 : _act_coefficient_a_2_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_2_T = act_op_sel_2 ? 32'h3e0c5859 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_2_T_1 = act_op_sel_1 ? 32'h3f000000 : _act_coefficient_b_2_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_2_T = act_op_sel_2 ? 32'h3f2c00da : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_2_T_1 = act_op_sel_1 ? 32'h3c9f42f6 : _act_coefficient_c_2_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_3_T = act_op_sel_2 ? 32'hba64a034 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_a_3_T_1 = act_op_sel_1 ? 32'hbc23b9f9 : _act_coefficient_a_3_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_3_T = act_op_sel_2 ? 32'h3c583b73 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_3_T_1 = act_op_sel_1 ? 32'h3f91554b : _act_coefficient_b_3_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_3_T = act_op_sel_2 ? 32'h3f731851 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_3_T_1 = act_op_sel_1 ? 32'hbeebfcc8 : _act_coefficient_c_3_T; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_b_4_T_1 = act_op_sel_1 ? 32'h3f800000 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_4_T = act_op_sel_2 ? 32'h3f800000 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_coefficient_c_4_T_1 = act_op_sel_1 ? 32'h0 : _act_coefficient_c_4_T; // @[Mux.scala 101:16]
  wire [31:0] _act_range_0_T_1 = act_op_sel_1 ? 32'hc1000000 : _act_coefficient_c_4_T; // @[Mux.scala 101:16]
  wire [31:0] _act_range_1_T = act_op_sel_2 ? 32'h40000000 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_range_1_T_1 = act_op_sel_1 ? 32'hc0000000 : _act_range_1_T; // @[Mux.scala 101:16]
  wire [31:0] _act_range_2_T = act_op_sel_2 ? 32'h40a00000 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_range_2_T_1 = act_op_sel_1 ? 32'h40000000 : _act_range_2_T; // @[Mux.scala 101:16]
  wire [31:0] _act_range_3_T = act_op_sel_2 ? 32'h41000000 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _act_range_3_T_1 = act_op_sel_1 ? 32'h41000000 : _act_range_3_T; // @[Mux.scala 101:16]
  wire [1:0] _act_func_prop_T = act_op_sel_2 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _act_func_prop_T_1 = act_op_sel_1 ? 2'h0 : _act_func_prop_T; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_a_0 = act_op_sel_0 ? 32'h0 : _act_coefficient_a_0_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_a_1 = act_op_sel_0 ? 32'h0 : _act_coefficient_a_1_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_a_2 = act_op_sel_0 ? 32'h0 : _act_coefficient_a_2_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_a_3 = act_op_sel_0 ? 32'h0 : _act_coefficient_a_3_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_b_0 = act_op_sel_0 ? 32'h0 : _act_coefficient_b_0_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_b_1 = act_op_sel_0 ? 32'h0 : _act_coefficient_b_1_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_b_2 = act_op_sel_0 ? 32'h0 : _act_coefficient_b_2_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_b_3 = act_op_sel_0 ? 32'h0 : _act_coefficient_b_3_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_b_4 = act_op_sel_0 ? 32'h0 : _act_coefficient_b_4_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_c_0 = act_op_sel_0 ? 32'h0 : _act_coefficient_c_0_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_c_1 = act_op_sel_0 ? 32'h0 : _act_coefficient_c_1_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_c_2 = act_op_sel_0 ? 32'h0 : _act_coefficient_c_2_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_c_3 = act_op_sel_0 ? 32'h0 : _act_coefficient_c_3_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_coefficient_c_4 = act_op_sel_0 ? 32'h0 : _act_coefficient_c_4_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_range_0 = act_op_sel_0 ? 32'h0 : _act_range_0_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_range_1 = act_op_sel_0 ? 32'h0 : _act_range_1_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_range_2 = act_op_sel_0 ? 32'h0 : _act_range_2_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_range_3 = act_op_sel_0 ? 32'h0 : _act_range_3_T_1; // @[Mux.scala 101:16]
  assign io_cfg_act_func_prop = act_op_sel_0 ? 2'h0 : _act_func_prop_T_1; // @[Mux.scala 101:16]
endmodule
module MuxOut(
  input         clock,
  input         reset,
  input  [31:0] io_i_data,
  input         io_cfg_act_en,
  input  [1:0]  io_act_func_prop,
  input  [31:0] io_cfg_coefficient_0,
  input  [31:0] io_cfg_coefficient_1,
  input  [31:0] io_cfg_coefficient_2,
  input  [31:0] io_cfg_coefficient_3,
  input  [31:0] io_cfg_coefficient_4,
  input  [31:0] io_x_range_0,
  input  [31:0] io_x_range_1,
  input  [31:0] io_x_range_2,
  input  [31:0] io_x_range_3,
  output [31:0] io_act_coefficient
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  act_prop = (io_act_func_prop == 2'h1 | io_act_func_prop == 2'h2) & io_i_data[31]; // @[act.scala 287:79]
  wire [31:0] _T_1 = {1'h0,io_i_data[30:0]}; // @[Cat.scala 33:92]
  wire [31:0] _T_2 = act_prop ? _T_1 : io_i_data; // @[act.scala 288:28]
  wire  _o_act_coefficient_T_9 = _T_2[31] ^ io_x_range_0[31] ? _T_2[31] : _T_2[30:0] < io_x_range_0[30:0] ^ _T_2[31]; // @[FP32.scala 48:8]
  wire  _o_act_coefficient_T_19 = _T_2[31] ^ io_x_range_1[31] ? _T_2[31] : _T_2[30:0] < io_x_range_1[30:0] ^ _T_2[31]; // @[FP32.scala 48:8]
  wire  _o_act_coefficient_T_29 = _T_2[31] ^ io_x_range_2[31] ? _T_2[31] : _T_2[30:0] < io_x_range_2[30:0] ^ _T_2[31]; // @[FP32.scala 48:8]
  wire  _o_act_coefficient_T_39 = _T_2[31] ^ io_x_range_3[31] ? _T_2[31] : _T_2[30:0] < io_x_range_3[30:0] ^ _T_2[31]; // @[FP32.scala 48:8]
  wire [31:0] _o_act_coefficient_T_40 = _o_act_coefficient_T_39 ? io_cfg_coefficient_3 : io_cfg_coefficient_4; // @[act.scala 299:62]
  wire [31:0] _o_act_coefficient_T_41 = _o_act_coefficient_T_29 ? io_cfg_coefficient_2 : _o_act_coefficient_T_40; // @[act.scala 299:16]
  reg [31:0] o_act_coefficient_t; // @[Reg.scala 35:20]
  assign io_act_coefficient = o_act_coefficient_t; // @[act.scala 304:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      o_act_coefficient_t <= 32'h0; // @[Reg.scala 35:20]
    end else if (io_cfg_act_en) begin // @[Reg.scala 36:18]
      if (_o_act_coefficient_T_9) begin // @[act.scala 293:32]
        o_act_coefficient_t <= io_cfg_coefficient_0;
      end else if (_o_act_coefficient_T_19) begin // @[act.scala 296:12]
        o_act_coefficient_t <= io_cfg_coefficient_1;
      end else begin
        o_act_coefficient_t <= _o_act_coefficient_T_41;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  o_act_coefficient_t = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module activationFuncDataCell(
  input         clock,
  input         reset,
  input  [31:0] io_i_data,
  input  [31:0] io_cfg_act_coefficient_a_0,
  input  [31:0] io_cfg_act_coefficient_a_1,
  input  [31:0] io_cfg_act_coefficient_a_2,
  input  [31:0] io_cfg_act_coefficient_a_3,
  input  [31:0] io_cfg_act_coefficient_b_0,
  input  [31:0] io_cfg_act_coefficient_b_1,
  input  [31:0] io_cfg_act_coefficient_b_2,
  input  [31:0] io_cfg_act_coefficient_b_3,
  input  [31:0] io_cfg_act_coefficient_b_4,
  input  [31:0] io_cfg_act_coefficient_c_0,
  input  [31:0] io_cfg_act_coefficient_c_1,
  input  [31:0] io_cfg_act_coefficient_c_2,
  input  [31:0] io_cfg_act_coefficient_c_3,
  input  [31:0] io_cfg_act_coefficient_c_4,
  input  [31:0] io_cfg_act_range_0,
  input  [31:0] io_cfg_act_range_1,
  input  [31:0] io_cfg_act_range_2,
  input  [31:0] io_cfg_act_range_3,
  input  [1:0]  io_cfg_act_func_prop,
  input  [1:0]  io_cfg_act_op,
  input         io_cfg_act_en,
  output [31:0] io_o_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
`endif // RANDOMIZE_REG_INIT
  wire  MuxOut_clock; // @[act.scala 315:36]
  wire  MuxOut_reset; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_i_data; // @[act.scala 315:36]
  wire  MuxOut_io_cfg_act_en; // @[act.scala 315:36]
  wire [1:0] MuxOut_io_act_func_prop; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_cfg_coefficient_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_cfg_coefficient_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_cfg_coefficient_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_cfg_coefficient_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_cfg_coefficient_4; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_x_range_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_x_range_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_x_range_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_x_range_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_io_act_coefficient; // @[act.scala 315:36]
  wire  MuxOut_1_clock; // @[act.scala 315:36]
  wire  MuxOut_1_reset; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_i_data; // @[act.scala 315:36]
  wire  MuxOut_1_io_cfg_act_en; // @[act.scala 315:36]
  wire [1:0] MuxOut_1_io_act_func_prop; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_cfg_coefficient_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_cfg_coefficient_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_cfg_coefficient_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_cfg_coefficient_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_cfg_coefficient_4; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_x_range_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_x_range_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_x_range_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_x_range_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_1_io_act_coefficient; // @[act.scala 315:36]
  wire  MuxOut_2_clock; // @[act.scala 315:36]
  wire  MuxOut_2_reset; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_i_data; // @[act.scala 315:36]
  wire  MuxOut_2_io_cfg_act_en; // @[act.scala 315:36]
  wire [1:0] MuxOut_2_io_act_func_prop; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_cfg_coefficient_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_cfg_coefficient_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_cfg_coefficient_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_cfg_coefficient_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_cfg_coefficient_4; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_x_range_0; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_x_range_1; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_x_range_2; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_x_range_3; // @[act.scala 315:36]
  wire [31:0] MuxOut_2_io_act_coefficient; // @[act.scala 315:36]
  wire  x_x_muler_clock; // @[Arithmetic.scala 95:25]
  wire  x_x_muler_reset; // @[Arithmetic.scala 95:25]
  wire [31:0] x_x_muler_io_x; // @[Arithmetic.scala 95:25]
  wire [31:0] x_x_muler_io_y; // @[Arithmetic.scala 95:25]
  wire [31:0] x_x_muler_io_z; // @[Arithmetic.scala 95:25]
  wire  x_x_muler_io_valid_in; // @[Arithmetic.scala 95:25]
  wire  x_b_muler_clock; // @[Arithmetic.scala 95:25]
  wire  x_b_muler_reset; // @[Arithmetic.scala 95:25]
  wire [31:0] x_b_muler_io_x; // @[Arithmetic.scala 95:25]
  wire [31:0] x_b_muler_io_y; // @[Arithmetic.scala 95:25]
  wire [31:0] x_b_muler_io_z; // @[Arithmetic.scala 95:25]
  wire  x_b_muler_io_valid_in; // @[Arithmetic.scala 95:25]
  wire  a_x_x_muler_clock; // @[Arithmetic.scala 95:25]
  wire  a_x_x_muler_reset; // @[Arithmetic.scala 95:25]
  wire [31:0] a_x_x_muler_io_x; // @[Arithmetic.scala 95:25]
  wire [31:0] a_x_x_muler_io_y; // @[Arithmetic.scala 95:25]
  wire [31:0] a_x_x_muler_io_z; // @[Arithmetic.scala 95:25]
  wire  a_x_x_muler_io_valid_in; // @[Arithmetic.scala 95:25]
  wire  x_b_and_c_adder_clock; // @[Arithmetic.scala 115:25]
  wire  x_b_and_c_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] x_b_and_c_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] x_b_and_c_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] x_b_and_c_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  x_b_and_c_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  axx_bx_c_adder_clock; // @[Arithmetic.scala 115:25]
  wire  axx_bx_c_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] axx_bx_c_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] axx_bx_c_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] axx_bx_c_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  axx_bx_c_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  io_o_data_adder_clock; // @[Arithmetic.scala 115:25]
  wire  io_o_data_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] io_o_data_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] io_o_data_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] io_o_data_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  io_o_data_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  reg [31:0] i_data_t; // @[act.scala 335:27]
  wire  _T_1 = io_cfg_act_func_prop == 2'h2; // @[act.scala 337:71]
  wire  _T_2 = io_cfg_act_func_prop == 2'h1 | io_cfg_act_func_prop == 2'h2; // @[act.scala 337:46]
  wire [31:0] _i_data_t_T_1 = {1'h0,io_i_data[30:0]}; // @[Cat.scala 33:92]
  reg [31:0] a_x_x_r; // @[Reg.scala 19:16]
  reg [31:0] x_b_and_c_r; // @[Reg.scala 19:16]
  reg [31:0] x_b_and_c_r_1; // @[Reg.scala 19:16]
  reg  i_sign_t_r; // @[Reg.scala 19:16]
  reg  i_sign_t_r_1; // @[Reg.scala 19:16]
  reg  i_sign_t_r_2; // @[Reg.scala 19:16]
  reg  i_sign_t_r_3; // @[Reg.scala 19:16]
  reg  i_sign_t_r_4; // @[Reg.scala 19:16]
  reg  i_sign_t_r_5; // @[Reg.scala 19:16]
  reg  i_sign_t_r_6; // @[Reg.scala 19:16]
  reg  i_sign_t_r_7; // @[Reg.scala 19:16]
  reg  i_sign_t_r_8; // @[Reg.scala 19:16]
  reg  i_sign_t_r_9; // @[Reg.scala 19:16]
  reg  i_sign_t_r_10; // @[Reg.scala 19:16]
  reg  i_sign_t_r_11; // @[Reg.scala 19:16]
  reg  i_sign_t; // @[Reg.scala 19:16]
  wire  o_data_prop = i_sign_t & _T_2; // @[act.scala 352:32]
  reg [31:0] axx_bx_c_r; // @[Reg.scala 19:16]
  wire [31:0] a_x_x_result_2_bits = a_x_x_muler_io_z; // @[Arithmetic.scala 124:22 125:17]
  reg [31:0] axx_bx_c_r_1; // @[Reg.scala 19:16]
  reg [31:0] axx_bx_c_r_2; // @[Reg.scala 19:16]
  reg [31:0] axx_bx_c_r_3; // @[Reg.scala 19:16]
  wire [31:0] axx_bx_c_bits = axx_bx_c_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire  _o_data_t_T_1 = ~axx_bx_c_bits[31]; // @[act.scala 361:42]
  wire [31:0] _o_data_t_T_3 = {_o_data_t_T_1,axx_bx_c_bits[30:0]}; // @[Cat.scala 33:92]
  reg  r; // @[Reg.scala 19:16]
  reg  r_1; // @[Reg.scala 19:16]
  reg  r_2; // @[Reg.scala 19:16]
  reg  r_3; // @[Reg.scala 19:16]
  reg  r_4; // @[Reg.scala 19:16]
  reg  r_5; // @[Reg.scala 19:16]
  reg  r_6; // @[Reg.scala 19:16]
  reg  r_7; // @[Reg.scala 19:16]
  reg  r_8; // @[Reg.scala 19:16]
  reg  r_9; // @[Reg.scala 19:16]
  reg  r_10; // @[Reg.scala 19:16]
  reg  r_11; // @[Reg.scala 19:16]
  reg  r_12; // @[Reg.scala 19:16]
  reg  r_13; // @[Reg.scala 19:16]
  reg  r_14; // @[Reg.scala 19:16]
  reg  r_15; // @[Reg.scala 19:16]
  reg  r_16; // @[Reg.scala 19:16]
  reg  r_17; // @[Reg.scala 19:16]
  reg [31:0] io_o_data_r; // @[Reg.scala 19:16]
  reg [31:0] io_o_data_r_1; // @[Reg.scala 19:16]
  reg [31:0] io_o_data_r_2; // @[Reg.scala 19:16]
  reg [31:0] io_o_data_r_3; // @[Reg.scala 19:16]
  reg [31:0] io_o_data_r_4; // @[Reg.scala 19:16]
  wire [31:0] io_o_data_result_2_bits = io_o_data_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] _GEN_45 = r_17 & _T_1 ? io_o_data_result_2_bits : io_o_data_r_4; // @[act.scala 366:129 367:19 369:19]
  MuxOut MuxOut ( // @[act.scala 315:36]
    .clock(MuxOut_clock),
    .reset(MuxOut_reset),
    .io_i_data(MuxOut_io_i_data),
    .io_cfg_act_en(MuxOut_io_cfg_act_en),
    .io_act_func_prop(MuxOut_io_act_func_prop),
    .io_cfg_coefficient_0(MuxOut_io_cfg_coefficient_0),
    .io_cfg_coefficient_1(MuxOut_io_cfg_coefficient_1),
    .io_cfg_coefficient_2(MuxOut_io_cfg_coefficient_2),
    .io_cfg_coefficient_3(MuxOut_io_cfg_coefficient_3),
    .io_cfg_coefficient_4(MuxOut_io_cfg_coefficient_4),
    .io_x_range_0(MuxOut_io_x_range_0),
    .io_x_range_1(MuxOut_io_x_range_1),
    .io_x_range_2(MuxOut_io_x_range_2),
    .io_x_range_3(MuxOut_io_x_range_3),
    .io_act_coefficient(MuxOut_io_act_coefficient)
  );
  MuxOut MuxOut_1 ( // @[act.scala 315:36]
    .clock(MuxOut_1_clock),
    .reset(MuxOut_1_reset),
    .io_i_data(MuxOut_1_io_i_data),
    .io_cfg_act_en(MuxOut_1_io_cfg_act_en),
    .io_act_func_prop(MuxOut_1_io_act_func_prop),
    .io_cfg_coefficient_0(MuxOut_1_io_cfg_coefficient_0),
    .io_cfg_coefficient_1(MuxOut_1_io_cfg_coefficient_1),
    .io_cfg_coefficient_2(MuxOut_1_io_cfg_coefficient_2),
    .io_cfg_coefficient_3(MuxOut_1_io_cfg_coefficient_3),
    .io_cfg_coefficient_4(MuxOut_1_io_cfg_coefficient_4),
    .io_x_range_0(MuxOut_1_io_x_range_0),
    .io_x_range_1(MuxOut_1_io_x_range_1),
    .io_x_range_2(MuxOut_1_io_x_range_2),
    .io_x_range_3(MuxOut_1_io_x_range_3),
    .io_act_coefficient(MuxOut_1_io_act_coefficient)
  );
  MuxOut MuxOut_2 ( // @[act.scala 315:36]
    .clock(MuxOut_2_clock),
    .reset(MuxOut_2_reset),
    .io_i_data(MuxOut_2_io_i_data),
    .io_cfg_act_en(MuxOut_2_io_cfg_act_en),
    .io_act_func_prop(MuxOut_2_io_act_func_prop),
    .io_cfg_coefficient_0(MuxOut_2_io_cfg_coefficient_0),
    .io_cfg_coefficient_1(MuxOut_2_io_cfg_coefficient_1),
    .io_cfg_coefficient_2(MuxOut_2_io_cfg_coefficient_2),
    .io_cfg_coefficient_3(MuxOut_2_io_cfg_coefficient_3),
    .io_cfg_coefficient_4(MuxOut_2_io_cfg_coefficient_4),
    .io_x_range_0(MuxOut_2_io_x_range_0),
    .io_x_range_1(MuxOut_2_io_x_range_1),
    .io_x_range_2(MuxOut_2_io_x_range_2),
    .io_x_range_3(MuxOut_2_io_x_range_3),
    .io_act_coefficient(MuxOut_2_io_act_coefficient)
  );
  FP32_Mult x_x_muler ( // @[Arithmetic.scala 95:25]
    .clock(x_x_muler_clock),
    .reset(x_x_muler_reset),
    .io_x(x_x_muler_io_x),
    .io_y(x_x_muler_io_y),
    .io_z(x_x_muler_io_z),
    .io_valid_in(x_x_muler_io_valid_in)
  );
  FP32_Mult x_b_muler ( // @[Arithmetic.scala 95:25]
    .clock(x_b_muler_clock),
    .reset(x_b_muler_reset),
    .io_x(x_b_muler_io_x),
    .io_y(x_b_muler_io_y),
    .io_z(x_b_muler_io_z),
    .io_valid_in(x_b_muler_io_valid_in)
  );
  FP32_Mult a_x_x_muler ( // @[Arithmetic.scala 95:25]
    .clock(a_x_x_muler_clock),
    .reset(a_x_x_muler_reset),
    .io_x(a_x_x_muler_io_x),
    .io_y(a_x_x_muler_io_y),
    .io_z(a_x_x_muler_io_z),
    .io_valid_in(a_x_x_muler_io_valid_in)
  );
  FP32_Adder x_b_and_c_adder ( // @[Arithmetic.scala 115:25]
    .clock(x_b_and_c_adder_clock),
    .reset(x_b_and_c_adder_reset),
    .io_x(x_b_and_c_adder_io_x),
    .io_y(x_b_and_c_adder_io_y),
    .io_z(x_b_and_c_adder_io_z),
    .io_valid_in(x_b_and_c_adder_io_valid_in)
  );
  FP32_Adder axx_bx_c_adder ( // @[Arithmetic.scala 115:25]
    .clock(axx_bx_c_adder_clock),
    .reset(axx_bx_c_adder_reset),
    .io_x(axx_bx_c_adder_io_x),
    .io_y(axx_bx_c_adder_io_y),
    .io_z(axx_bx_c_adder_io_z),
    .io_valid_in(axx_bx_c_adder_io_valid_in)
  );
  FP32_Adder io_o_data_adder ( // @[Arithmetic.scala 115:25]
    .clock(io_o_data_adder_clock),
    .reset(io_o_data_adder_reset),
    .io_x(io_o_data_adder_io_x),
    .io_y(io_o_data_adder_io_y),
    .io_z(io_o_data_adder_io_z),
    .io_valid_in(io_o_data_adder_io_valid_in)
  );
  assign io_o_data = io_cfg_act_op == 2'h0 ? io_i_data : _GEN_45; // @[act.scala 364:33 365:19]
  assign MuxOut_clock = clock;
  assign MuxOut_reset = reset;
  assign MuxOut_io_i_data = io_i_data; // @[act.scala 318:33]
  assign MuxOut_io_cfg_act_en = io_cfg_act_en; // @[act.scala 319:33]
  assign MuxOut_io_act_func_prop = io_cfg_act_func_prop; // @[act.scala 320:33]
  assign MuxOut_io_cfg_coefficient_0 = io_cfg_act_coefficient_a_0; // @[act.scala 323:31]
  assign MuxOut_io_cfg_coefficient_1 = io_cfg_act_coefficient_a_1; // @[act.scala 323:31]
  assign MuxOut_io_cfg_coefficient_2 = io_cfg_act_coefficient_a_2; // @[act.scala 323:31]
  assign MuxOut_io_cfg_coefficient_3 = io_cfg_act_coefficient_a_3; // @[act.scala 323:31]
  assign MuxOut_io_cfg_coefficient_4 = 32'h0; // @[act.scala 323:31]
  assign MuxOut_io_x_range_0 = io_cfg_act_range_0; // @[act.scala 321:33]
  assign MuxOut_io_x_range_1 = io_cfg_act_range_1; // @[act.scala 321:33]
  assign MuxOut_io_x_range_2 = io_cfg_act_range_2; // @[act.scala 321:33]
  assign MuxOut_io_x_range_3 = io_cfg_act_range_3; // @[act.scala 321:33]
  assign MuxOut_1_clock = clock;
  assign MuxOut_1_reset = reset;
  assign MuxOut_1_io_i_data = io_i_data; // @[act.scala 318:33]
  assign MuxOut_1_io_cfg_act_en = io_cfg_act_en; // @[act.scala 319:33]
  assign MuxOut_1_io_act_func_prop = io_cfg_act_func_prop; // @[act.scala 320:33]
  assign MuxOut_1_io_cfg_coefficient_0 = io_cfg_act_coefficient_b_0; // @[act.scala 324:31]
  assign MuxOut_1_io_cfg_coefficient_1 = io_cfg_act_coefficient_b_1; // @[act.scala 324:31]
  assign MuxOut_1_io_cfg_coefficient_2 = io_cfg_act_coefficient_b_2; // @[act.scala 324:31]
  assign MuxOut_1_io_cfg_coefficient_3 = io_cfg_act_coefficient_b_3; // @[act.scala 324:31]
  assign MuxOut_1_io_cfg_coefficient_4 = io_cfg_act_coefficient_b_4; // @[act.scala 324:31]
  assign MuxOut_1_io_x_range_0 = io_cfg_act_range_0; // @[act.scala 321:33]
  assign MuxOut_1_io_x_range_1 = io_cfg_act_range_1; // @[act.scala 321:33]
  assign MuxOut_1_io_x_range_2 = io_cfg_act_range_2; // @[act.scala 321:33]
  assign MuxOut_1_io_x_range_3 = io_cfg_act_range_3; // @[act.scala 321:33]
  assign MuxOut_2_clock = clock;
  assign MuxOut_2_reset = reset;
  assign MuxOut_2_io_i_data = io_i_data; // @[act.scala 318:33]
  assign MuxOut_2_io_cfg_act_en = io_cfg_act_en; // @[act.scala 319:33]
  assign MuxOut_2_io_act_func_prop = io_cfg_act_func_prop; // @[act.scala 320:33]
  assign MuxOut_2_io_cfg_coefficient_0 = io_cfg_act_coefficient_c_0; // @[act.scala 325:31]
  assign MuxOut_2_io_cfg_coefficient_1 = io_cfg_act_coefficient_c_1; // @[act.scala 325:31]
  assign MuxOut_2_io_cfg_coefficient_2 = io_cfg_act_coefficient_c_2; // @[act.scala 325:31]
  assign MuxOut_2_io_cfg_coefficient_3 = io_cfg_act_coefficient_c_3; // @[act.scala 325:31]
  assign MuxOut_2_io_cfg_coefficient_4 = io_cfg_act_coefficient_c_4; // @[act.scala 325:31]
  assign MuxOut_2_io_x_range_0 = io_cfg_act_range_0; // @[act.scala 321:33]
  assign MuxOut_2_io_x_range_1 = io_cfg_act_range_1; // @[act.scala 321:33]
  assign MuxOut_2_io_x_range_2 = io_cfg_act_range_2; // @[act.scala 321:33]
  assign MuxOut_2_io_x_range_3 = io_cfg_act_range_3; // @[act.scala 321:33]
  assign x_x_muler_clock = clock;
  assign x_x_muler_reset = reset;
  assign x_x_muler_io_x = io_i_data; // @[Arithmetic.scala 124:22 125:17]
  assign x_x_muler_io_y = io_i_data; // @[Arithmetic.scala 124:22 125:17]
  assign x_x_muler_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 98:25]
  assign x_b_muler_clock = clock;
  assign x_b_muler_reset = reset;
  assign x_b_muler_io_x = i_data_t; // @[Arithmetic.scala 124:22 125:17]
  assign x_b_muler_io_y = MuxOut_1_io_act_coefficient; // @[Arithmetic.scala 124:22 125:17]
  assign x_b_muler_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 98:25]
  assign a_x_x_muler_clock = clock;
  assign a_x_x_muler_reset = reset;
  assign a_x_x_muler_io_x = a_x_x_r; // @[Arithmetic.scala 124:22 125:17]
  assign a_x_x_muler_io_y = x_x_muler_io_z; // @[Arithmetic.scala 124:22 125:17]
  assign a_x_x_muler_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 98:25]
  assign x_b_and_c_adder_clock = clock;
  assign x_b_and_c_adder_reset = reset;
  assign x_b_and_c_adder_io_x = x_b_and_c_r_1; // @[Arithmetic.scala 124:22 125:17]
  assign x_b_and_c_adder_io_y = x_b_muler_io_z; // @[Arithmetic.scala 124:22 125:17]
  assign x_b_and_c_adder_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 118:25]
  assign axx_bx_c_adder_clock = clock;
  assign axx_bx_c_adder_reset = reset;
  assign axx_bx_c_adder_io_x = axx_bx_c_r_3; // @[Arithmetic.scala 124:22 125:17]
  assign axx_bx_c_adder_io_y = x_b_and_c_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  assign axx_bx_c_adder_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 118:25]
  assign io_o_data_adder_clock = clock;
  assign io_o_data_adder_reset = reset;
  assign io_o_data_adder_io_x = o_data_prop ? _o_data_t_T_3 : axx_bx_c_bits; // @[act.scala 361:24]
  assign io_o_data_adder_io_y = 32'h3f800000; // @[Arithmetic.scala 124:22 125:17]
  assign io_o_data_adder_io_valid_in = io_cfg_act_en; // @[Arithmetic.scala 118:25]
  always @(posedge clock) begin
    if (reset) begin // @[act.scala 335:27]
      i_data_t <= 32'h0; // @[act.scala 335:27]
    end else if (io_cfg_act_en) begin // @[act.scala 336:24]
      if ((io_cfg_act_func_prop == 2'h1 | io_cfg_act_func_prop == 2'h2) & io_i_data[31]) begin // @[act.scala 337:108]
        i_data_t <= _i_data_t_T_1; // @[act.scala 338:22]
      end else begin
        i_data_t <= io_i_data; // @[act.scala 340:22]
      end
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      a_x_x_r <= MuxOut_io_act_coefficient; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      x_b_and_c_r <= MuxOut_2_io_act_coefficient; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      x_b_and_c_r_1 <= x_b_and_c_r; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r <= io_i_data[31]; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_1 <= i_sign_t_r; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_2 <= i_sign_t_r_1; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_3 <= i_sign_t_r_2; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_4 <= i_sign_t_r_3; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_5 <= i_sign_t_r_4; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_6 <= i_sign_t_r_5; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_7 <= i_sign_t_r_6; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_8 <= i_sign_t_r_7; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_9 <= i_sign_t_r_8; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_10 <= i_sign_t_r_9; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t_r_11 <= i_sign_t_r_10; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      i_sign_t <= i_sign_t_r_11; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      axx_bx_c_r <= a_x_x_result_2_bits; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      axx_bx_c_r_1 <= axx_bx_c_r; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      axx_bx_c_r_2 <= axx_bx_c_r_1; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      axx_bx_c_r_3 <= axx_bx_c_r_2; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r <= io_i_data[31]; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_1 <= r; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_2 <= r_1; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_3 <= r_2; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_4 <= r_3; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_5 <= r_4; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_6 <= r_5; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_7 <= r_6; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_8 <= r_7; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_9 <= r_8; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_10 <= r_9; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_11 <= r_10; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_12 <= r_11; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_13 <= r_12; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_14 <= r_13; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_15 <= r_14; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_16 <= r_15; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      r_17 <= r_16; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      if (o_data_prop) begin // @[act.scala 361:24]
        io_o_data_r <= _o_data_t_T_3;
      end else begin
        io_o_data_r <= axx_bx_c_bits;
      end
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      io_o_data_r_1 <= io_o_data_r; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      io_o_data_r_2 <= io_o_data_r_1; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      io_o_data_r_3 <= io_o_data_r_2; // @[Reg.scala 20:22]
    end
    if (io_cfg_act_en) begin // @[Reg.scala 20:18]
      io_o_data_r_4 <= io_o_data_r_3; // @[Reg.scala 20:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  i_data_t = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  a_x_x_r = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_b_and_c_r = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_b_and_c_r_1 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  i_sign_t_r = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  i_sign_t_r_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  i_sign_t_r_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  i_sign_t_r_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  i_sign_t_r_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  i_sign_t_r_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  i_sign_t_r_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  i_sign_t_r_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  i_sign_t_r_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  i_sign_t_r_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  i_sign_t_r_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  i_sign_t_r_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  i_sign_t = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  axx_bx_c_r = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  axx_bx_c_r_1 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  axx_bx_c_r_2 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  axx_bx_c_r_3 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  r = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  r_1 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  r_2 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  r_3 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  r_4 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  r_5 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  r_6 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  r_7 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  r_8 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  r_9 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  r_10 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  r_11 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  r_12 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  r_13 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  r_14 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  r_15 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  r_16 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  r_17 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  io_o_data_r = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  io_o_data_r_1 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  io_o_data_r_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  io_o_data_r_3 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  io_o_data_r_4 = _RAND_43[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module activationFunc(
  input         clock,
  input         reset,
  input  [31:0] io_cfg_act_coefficient_a_0,
  input  [31:0] io_cfg_act_coefficient_a_1,
  input  [31:0] io_cfg_act_coefficient_a_2,
  input  [31:0] io_cfg_act_coefficient_a_3,
  input  [31:0] io_cfg_act_coefficient_b_0,
  input  [31:0] io_cfg_act_coefficient_b_1,
  input  [31:0] io_cfg_act_coefficient_b_2,
  input  [31:0] io_cfg_act_coefficient_b_3,
  input  [31:0] io_cfg_act_coefficient_b_4,
  input  [31:0] io_cfg_act_coefficient_c_0,
  input  [31:0] io_cfg_act_coefficient_c_1,
  input  [31:0] io_cfg_act_coefficient_c_2,
  input  [31:0] io_cfg_act_coefficient_c_3,
  input  [31:0] io_cfg_act_coefficient_c_4,
  input  [31:0] io_cfg_act_range_0,
  input  [31:0] io_cfg_act_range_1,
  input  [31:0] io_cfg_act_range_2,
  input  [31:0] io_cfg_act_range_3,
  input  [1:0]  io_cfg_act_func_prop,
  input  [1:0]  io_cfg_act_op,
  input         io_cfg_act_en,
  input  [31:0] io_i_data_data_0,
  input  [31:0] io_i_data_data_1,
  input  [31:0] io_i_data_data_2,
  input  [31:0] io_i_data_data_3,
  input  [31:0] io_i_data_data_4,
  input  [31:0] io_i_data_data_5,
  input  [31:0] io_i_data_data_6,
  input  [31:0] io_i_data_data_7,
  output [31:0] io_o_data_data_0,
  output [31:0] io_o_data_data_1,
  output [31:0] io_o_data_data_2,
  output [31:0] io_o_data_data_3,
  output [31:0] io_o_data_data_4,
  output [31:0] io_o_data_data_5,
  output [31:0] io_o_data_data_6,
  output [31:0] io_o_data_data_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  wire  activationFuncDataCell_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_1_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_1_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_1_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_1_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_1_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_1_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_2_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_2_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_2_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_2_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_2_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_2_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_3_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_3_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_3_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_3_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_3_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_3_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_4_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_4_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_4_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_4_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_4_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_4_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_5_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_5_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_5_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_5_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_5_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_5_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_6_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_6_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_6_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_6_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_6_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_6_io_o_data; // @[act.scala 242:57]
  wire  activationFuncDataCell_7_clock; // @[act.scala 242:57]
  wire  activationFuncDataCell_7_reset; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_i_data; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_a_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_a_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_a_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_a_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_b_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_b_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_b_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_b_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_b_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_c_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_c_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_c_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_c_3; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_coefficient_c_4; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_range_0; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_range_1; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_range_2; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_cfg_act_range_3; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_7_io_cfg_act_func_prop; // @[act.scala 242:57]
  wire [1:0] activationFuncDataCell_7_io_cfg_act_op; // @[act.scala 242:57]
  wire  activationFuncDataCell_7_io_cfg_act_en; // @[act.scala 242:57]
  wire [31:0] activationFuncDataCell_7_io_o_data; // @[act.scala 242:57]
  reg  cfg_REG; // @[utils.scala 28:16]
  wire  _cfg_T = cfg_REG ^ io_cfg_act_en; // @[utils.scala 28:26]
  reg [31:0] cfg_act_coefficient_a_0; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_a_1; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_a_2; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_a_3; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_b_0; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_b_1; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_b_2; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_b_3; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_b_4; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_c_0; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_c_1; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_c_2; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_c_3; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_coefficient_c_4; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_range_0; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_range_1; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_range_2; // @[Reg.scala 35:20]
  reg [31:0] cfg_act_range_3; // @[Reg.scala 35:20]
  reg [1:0] cfg_act_func_prop; // @[Reg.scala 35:20]
  reg [1:0] cfg_act_op; // @[Reg.scala 35:20]
  reg  cfg_act_en; // @[Reg.scala 35:20]
  activationFuncDataCell activationFuncDataCell ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_clock),
    .reset(activationFuncDataCell_reset),
    .io_i_data(activationFuncDataCell_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_1 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_1_clock),
    .reset(activationFuncDataCell_1_reset),
    .io_i_data(activationFuncDataCell_1_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_1_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_1_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_1_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_1_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_1_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_1_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_1_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_1_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_1_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_1_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_1_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_1_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_1_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_1_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_1_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_1_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_1_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_1_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_1_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_1_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_1_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_1_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_2 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_2_clock),
    .reset(activationFuncDataCell_2_reset),
    .io_i_data(activationFuncDataCell_2_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_2_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_2_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_2_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_2_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_2_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_2_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_2_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_2_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_2_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_2_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_2_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_2_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_2_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_2_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_2_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_2_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_2_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_2_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_2_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_2_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_2_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_2_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_3 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_3_clock),
    .reset(activationFuncDataCell_3_reset),
    .io_i_data(activationFuncDataCell_3_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_3_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_3_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_3_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_3_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_3_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_3_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_3_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_3_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_3_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_3_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_3_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_3_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_3_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_3_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_3_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_3_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_3_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_3_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_3_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_3_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_3_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_3_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_4 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_4_clock),
    .reset(activationFuncDataCell_4_reset),
    .io_i_data(activationFuncDataCell_4_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_4_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_4_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_4_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_4_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_4_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_4_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_4_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_4_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_4_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_4_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_4_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_4_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_4_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_4_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_4_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_4_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_4_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_4_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_4_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_4_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_4_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_4_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_5 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_5_clock),
    .reset(activationFuncDataCell_5_reset),
    .io_i_data(activationFuncDataCell_5_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_5_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_5_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_5_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_5_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_5_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_5_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_5_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_5_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_5_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_5_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_5_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_5_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_5_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_5_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_5_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_5_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_5_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_5_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_5_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_5_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_5_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_5_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_6 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_6_clock),
    .reset(activationFuncDataCell_6_reset),
    .io_i_data(activationFuncDataCell_6_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_6_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_6_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_6_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_6_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_6_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_6_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_6_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_6_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_6_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_6_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_6_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_6_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_6_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_6_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_6_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_6_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_6_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_6_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_6_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_6_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_6_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_6_io_o_data)
  );
  activationFuncDataCell activationFuncDataCell_7 ( // @[act.scala 242:57]
    .clock(activationFuncDataCell_7_clock),
    .reset(activationFuncDataCell_7_reset),
    .io_i_data(activationFuncDataCell_7_io_i_data),
    .io_cfg_act_coefficient_a_0(activationFuncDataCell_7_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(activationFuncDataCell_7_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(activationFuncDataCell_7_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(activationFuncDataCell_7_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(activationFuncDataCell_7_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(activationFuncDataCell_7_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(activationFuncDataCell_7_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(activationFuncDataCell_7_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(activationFuncDataCell_7_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(activationFuncDataCell_7_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(activationFuncDataCell_7_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(activationFuncDataCell_7_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(activationFuncDataCell_7_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(activationFuncDataCell_7_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(activationFuncDataCell_7_io_cfg_act_range_0),
    .io_cfg_act_range_1(activationFuncDataCell_7_io_cfg_act_range_1),
    .io_cfg_act_range_2(activationFuncDataCell_7_io_cfg_act_range_2),
    .io_cfg_act_range_3(activationFuncDataCell_7_io_cfg_act_range_3),
    .io_cfg_act_func_prop(activationFuncDataCell_7_io_cfg_act_func_prop),
    .io_cfg_act_op(activationFuncDataCell_7_io_cfg_act_op),
    .io_cfg_act_en(activationFuncDataCell_7_io_cfg_act_en),
    .io_o_data(activationFuncDataCell_7_io_o_data)
  );
  assign io_o_data_data_0 = activationFuncDataCell_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_1 = activationFuncDataCell_1_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_2 = activationFuncDataCell_2_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_3 = activationFuncDataCell_3_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_4 = activationFuncDataCell_4_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_5 = activationFuncDataCell_5_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_6 = activationFuncDataCell_6_io_o_data; // @[act.scala 252:42]
  assign io_o_data_data_7 = activationFuncDataCell_7_io_o_data; // @[act.scala 252:42]
  assign activationFuncDataCell_clock = clock;
  assign activationFuncDataCell_reset = reset;
  assign activationFuncDataCell_io_i_data = io_i_data_data_0; // @[act.scala 250:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_1_clock = clock;
  assign activationFuncDataCell_1_reset = reset;
  assign activationFuncDataCell_1_io_i_data = io_i_data_data_1; // @[act.scala 250:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_1_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_2_clock = clock;
  assign activationFuncDataCell_2_reset = reset;
  assign activationFuncDataCell_2_io_i_data = io_i_data_data_2; // @[act.scala 250:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_2_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_3_clock = clock;
  assign activationFuncDataCell_3_reset = reset;
  assign activationFuncDataCell_3_io_i_data = io_i_data_data_3; // @[act.scala 250:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_3_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_4_clock = clock;
  assign activationFuncDataCell_4_reset = reset;
  assign activationFuncDataCell_4_io_i_data = io_i_data_data_4; // @[act.scala 250:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_4_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_5_clock = clock;
  assign activationFuncDataCell_5_reset = reset;
  assign activationFuncDataCell_5_io_i_data = io_i_data_data_5; // @[act.scala 250:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_5_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_6_clock = clock;
  assign activationFuncDataCell_6_reset = reset;
  assign activationFuncDataCell_6_io_i_data = io_i_data_data_6; // @[act.scala 250:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_6_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  assign activationFuncDataCell_7_clock = clock;
  assign activationFuncDataCell_7_reset = reset;
  assign activationFuncDataCell_7_io_i_data = io_i_data_data_7; // @[act.scala 250:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_a_0 = cfg_act_coefficient_a_0; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_a_1 = cfg_act_coefficient_a_1; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_a_2 = cfg_act_coefficient_a_2; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_a_3 = cfg_act_coefficient_a_3; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_b_0 = cfg_act_coefficient_b_0; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_b_1 = cfg_act_coefficient_b_1; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_b_2 = cfg_act_coefficient_b_2; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_b_3 = cfg_act_coefficient_b_3; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_b_4 = cfg_act_coefficient_b_4; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_c_0 = cfg_act_coefficient_c_0; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_c_1 = cfg_act_coefficient_c_1; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_c_2 = cfg_act_coefficient_c_2; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_c_3 = cfg_act_coefficient_c_3; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_coefficient_c_4 = cfg_act_coefficient_c_4; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_range_0 = cfg_act_range_0; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_range_1 = cfg_act_range_1; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_range_2 = cfg_act_range_2; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_range_3 = cfg_act_range_3; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_func_prop = cfg_act_func_prop; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_op = cfg_act_op; // @[act.scala 251:42]
  assign activationFuncDataCell_7_io_cfg_act_en = cfg_act_en; // @[act.scala 251:42]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 28:16]
      cfg_REG <= 1'h0; // @[utils.scala 28:16]
    end else begin
      cfg_REG <= io_cfg_act_en; // @[utils.scala 28:16]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_a_0 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_a_0 <= io_cfg_act_coefficient_a_0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_a_1 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_a_1 <= io_cfg_act_coefficient_a_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_a_2 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_a_2 <= io_cfg_act_coefficient_a_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_a_3 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_a_3 <= io_cfg_act_coefficient_a_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_b_0 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_b_0 <= io_cfg_act_coefficient_b_0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_b_1 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_b_1 <= io_cfg_act_coefficient_b_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_b_2 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_b_2 <= io_cfg_act_coefficient_b_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_b_3 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_b_3 <= io_cfg_act_coefficient_b_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_b_4 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_b_4 <= io_cfg_act_coefficient_b_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_c_0 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_c_0 <= io_cfg_act_coefficient_c_0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_c_1 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_c_1 <= io_cfg_act_coefficient_c_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_c_2 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_c_2 <= io_cfg_act_coefficient_c_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_c_3 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_c_3 <= io_cfg_act_coefficient_c_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_coefficient_c_4 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_coefficient_c_4 <= io_cfg_act_coefficient_c_4; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_range_0 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_range_0 <= io_cfg_act_range_0; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_range_1 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_range_1 <= io_cfg_act_range_1; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_range_2 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_range_2 <= io_cfg_act_range_2; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_range_3 <= 32'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_range_3 <= io_cfg_act_range_3; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_func_prop <= 2'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_func_prop <= io_cfg_act_func_prop; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_op <= 2'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_op <= io_cfg_act_op; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      cfg_act_en <= 1'h0; // @[Reg.scala 35:20]
    end else if (_cfg_T) begin // @[Reg.scala 36:18]
      cfg_act_en <= io_cfg_act_en; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cfg_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cfg_act_coefficient_a_0 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  cfg_act_coefficient_a_1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cfg_act_coefficient_a_2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cfg_act_coefficient_a_3 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cfg_act_coefficient_b_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cfg_act_coefficient_b_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  cfg_act_coefficient_b_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  cfg_act_coefficient_b_3 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  cfg_act_coefficient_b_4 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cfg_act_coefficient_c_0 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  cfg_act_coefficient_c_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  cfg_act_coefficient_c_2 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  cfg_act_coefficient_c_3 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  cfg_act_coefficient_c_4 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  cfg_act_range_0 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  cfg_act_range_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  cfg_act_range_2 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  cfg_act_range_3 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  cfg_act_func_prop = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  cfg_act_op = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  cfg_act_en = _RAND_21[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module alu_act(
  input         clock,
  input         reset,
  input  [1:0]  io_act_op,
  input         io_act_en,
  input  [31:0] io_i_data_data_0,
  input  [31:0] io_i_data_data_1,
  input  [31:0] io_i_data_data_2,
  input  [31:0] io_i_data_data_3,
  input  [31:0] io_i_data_data_4,
  input  [31:0] io_i_data_data_5,
  input  [31:0] io_i_data_data_6,
  input  [31:0] io_i_data_data_7,
  output [31:0] io_o_data_data_0,
  output [31:0] io_o_data_data_1,
  output [31:0] io_o_data_data_2,
  output [31:0] io_o_data_data_3,
  output [31:0] io_o_data_data_4,
  output [31:0] io_o_data_data_5,
  output [31:0] io_o_data_data_6,
  output [31:0] io_o_data_data_7
);
  wire [1:0] alu_act_param_select_io_act_op; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_a_0; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_a_1; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_a_2; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_a_3; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_b_0; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_b_1; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_b_2; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_b_3; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_b_4; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_c_0; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_c_1; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_c_2; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_c_3; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_coefficient_c_4; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_range_0; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_range_1; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_range_2; // @[act.scala 122:38]
  wire [31:0] alu_act_param_select_io_cfg_act_range_3; // @[act.scala 122:38]
  wire [1:0] alu_act_param_select_io_cfg_act_func_prop; // @[act.scala 122:38]
  wire  actfunc_clock; // @[act.scala 135:25]
  wire  actfunc_reset; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_a_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_a_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_a_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_a_3; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_b_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_b_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_b_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_b_3; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_b_4; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_c_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_c_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_c_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_c_3; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_coefficient_c_4; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_range_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_range_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_range_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_cfg_act_range_3; // @[act.scala 135:25]
  wire [1:0] actfunc_io_cfg_act_func_prop; // @[act.scala 135:25]
  wire [1:0] actfunc_io_cfg_act_op; // @[act.scala 135:25]
  wire  actfunc_io_cfg_act_en; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_3; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_4; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_5; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_6; // @[act.scala 135:25]
  wire [31:0] actfunc_io_i_data_data_7; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_0; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_1; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_2; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_3; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_4; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_5; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_6; // @[act.scala 135:25]
  wire [31:0] actfunc_io_o_data_data_7; // @[act.scala 135:25]
  alu_act_param_select alu_act_param_select ( // @[act.scala 122:38]
    .io_act_op(alu_act_param_select_io_act_op),
    .io_cfg_act_coefficient_a_0(alu_act_param_select_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(alu_act_param_select_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(alu_act_param_select_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(alu_act_param_select_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(alu_act_param_select_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(alu_act_param_select_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(alu_act_param_select_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(alu_act_param_select_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(alu_act_param_select_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(alu_act_param_select_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(alu_act_param_select_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(alu_act_param_select_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(alu_act_param_select_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(alu_act_param_select_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(alu_act_param_select_io_cfg_act_range_0),
    .io_cfg_act_range_1(alu_act_param_select_io_cfg_act_range_1),
    .io_cfg_act_range_2(alu_act_param_select_io_cfg_act_range_2),
    .io_cfg_act_range_3(alu_act_param_select_io_cfg_act_range_3),
    .io_cfg_act_func_prop(alu_act_param_select_io_cfg_act_func_prop)
  );
  activationFunc actfunc ( // @[act.scala 135:25]
    .clock(actfunc_clock),
    .reset(actfunc_reset),
    .io_cfg_act_coefficient_a_0(actfunc_io_cfg_act_coefficient_a_0),
    .io_cfg_act_coefficient_a_1(actfunc_io_cfg_act_coefficient_a_1),
    .io_cfg_act_coefficient_a_2(actfunc_io_cfg_act_coefficient_a_2),
    .io_cfg_act_coefficient_a_3(actfunc_io_cfg_act_coefficient_a_3),
    .io_cfg_act_coefficient_b_0(actfunc_io_cfg_act_coefficient_b_0),
    .io_cfg_act_coefficient_b_1(actfunc_io_cfg_act_coefficient_b_1),
    .io_cfg_act_coefficient_b_2(actfunc_io_cfg_act_coefficient_b_2),
    .io_cfg_act_coefficient_b_3(actfunc_io_cfg_act_coefficient_b_3),
    .io_cfg_act_coefficient_b_4(actfunc_io_cfg_act_coefficient_b_4),
    .io_cfg_act_coefficient_c_0(actfunc_io_cfg_act_coefficient_c_0),
    .io_cfg_act_coefficient_c_1(actfunc_io_cfg_act_coefficient_c_1),
    .io_cfg_act_coefficient_c_2(actfunc_io_cfg_act_coefficient_c_2),
    .io_cfg_act_coefficient_c_3(actfunc_io_cfg_act_coefficient_c_3),
    .io_cfg_act_coefficient_c_4(actfunc_io_cfg_act_coefficient_c_4),
    .io_cfg_act_range_0(actfunc_io_cfg_act_range_0),
    .io_cfg_act_range_1(actfunc_io_cfg_act_range_1),
    .io_cfg_act_range_2(actfunc_io_cfg_act_range_2),
    .io_cfg_act_range_3(actfunc_io_cfg_act_range_3),
    .io_cfg_act_func_prop(actfunc_io_cfg_act_func_prop),
    .io_cfg_act_op(actfunc_io_cfg_act_op),
    .io_cfg_act_en(actfunc_io_cfg_act_en),
    .io_i_data_data_0(actfunc_io_i_data_data_0),
    .io_i_data_data_1(actfunc_io_i_data_data_1),
    .io_i_data_data_2(actfunc_io_i_data_data_2),
    .io_i_data_data_3(actfunc_io_i_data_data_3),
    .io_i_data_data_4(actfunc_io_i_data_data_4),
    .io_i_data_data_5(actfunc_io_i_data_data_5),
    .io_i_data_data_6(actfunc_io_i_data_data_6),
    .io_i_data_data_7(actfunc_io_i_data_data_7),
    .io_o_data_data_0(actfunc_io_o_data_data_0),
    .io_o_data_data_1(actfunc_io_o_data_data_1),
    .io_o_data_data_2(actfunc_io_o_data_data_2),
    .io_o_data_data_3(actfunc_io_o_data_data_3),
    .io_o_data_data_4(actfunc_io_o_data_data_4),
    .io_o_data_data_5(actfunc_io_o_data_data_5),
    .io_o_data_data_6(actfunc_io_o_data_data_6),
    .io_o_data_data_7(actfunc_io_o_data_data_7)
  );
  assign io_o_data_data_0 = actfunc_io_o_data_data_0; // @[act.scala 138:15]
  assign io_o_data_data_1 = actfunc_io_o_data_data_1; // @[act.scala 138:15]
  assign io_o_data_data_2 = actfunc_io_o_data_data_2; // @[act.scala 138:15]
  assign io_o_data_data_3 = actfunc_io_o_data_data_3; // @[act.scala 138:15]
  assign io_o_data_data_4 = actfunc_io_o_data_data_4; // @[act.scala 138:15]
  assign io_o_data_data_5 = actfunc_io_o_data_data_5; // @[act.scala 138:15]
  assign io_o_data_data_6 = actfunc_io_o_data_data_6; // @[act.scala 138:15]
  assign io_o_data_data_7 = actfunc_io_o_data_data_7; // @[act.scala 138:15]
  assign alu_act_param_select_io_act_op = io_act_op; // @[act.scala 128:35]
  assign actfunc_clock = clock;
  assign actfunc_reset = reset;
  assign actfunc_io_cfg_act_coefficient_a_0 = alu_act_param_select_io_cfg_act_coefficient_a_0; // @[act.scala 124:19 130:27]
  assign actfunc_io_cfg_act_coefficient_a_1 = alu_act_param_select_io_cfg_act_coefficient_a_1; // @[act.scala 124:19 130:27]
  assign actfunc_io_cfg_act_coefficient_a_2 = alu_act_param_select_io_cfg_act_coefficient_a_2; // @[act.scala 124:19 130:27]
  assign actfunc_io_cfg_act_coefficient_a_3 = alu_act_param_select_io_cfg_act_coefficient_a_3; // @[act.scala 124:19 130:27]
  assign actfunc_io_cfg_act_coefficient_b_0 = alu_act_param_select_io_cfg_act_coefficient_b_0; // @[act.scala 124:19 131:27]
  assign actfunc_io_cfg_act_coefficient_b_1 = alu_act_param_select_io_cfg_act_coefficient_b_1; // @[act.scala 124:19 131:27]
  assign actfunc_io_cfg_act_coefficient_b_2 = alu_act_param_select_io_cfg_act_coefficient_b_2; // @[act.scala 124:19 131:27]
  assign actfunc_io_cfg_act_coefficient_b_3 = alu_act_param_select_io_cfg_act_coefficient_b_3; // @[act.scala 124:19 131:27]
  assign actfunc_io_cfg_act_coefficient_b_4 = alu_act_param_select_io_cfg_act_coefficient_b_4; // @[act.scala 124:19 131:27]
  assign actfunc_io_cfg_act_coefficient_c_0 = alu_act_param_select_io_cfg_act_coefficient_c_0; // @[act.scala 124:19 132:27]
  assign actfunc_io_cfg_act_coefficient_c_1 = alu_act_param_select_io_cfg_act_coefficient_c_1; // @[act.scala 124:19 132:27]
  assign actfunc_io_cfg_act_coefficient_c_2 = alu_act_param_select_io_cfg_act_coefficient_c_2; // @[act.scala 124:19 132:27]
  assign actfunc_io_cfg_act_coefficient_c_3 = alu_act_param_select_io_cfg_act_coefficient_c_3; // @[act.scala 124:19 132:27]
  assign actfunc_io_cfg_act_coefficient_c_4 = alu_act_param_select_io_cfg_act_coefficient_c_4; // @[act.scala 124:19 132:27]
  assign actfunc_io_cfg_act_range_0 = alu_act_param_select_io_cfg_act_range_0; // @[act.scala 124:19 129:19]
  assign actfunc_io_cfg_act_range_1 = alu_act_param_select_io_cfg_act_range_1; // @[act.scala 124:19 129:19]
  assign actfunc_io_cfg_act_range_2 = alu_act_param_select_io_cfg_act_range_2; // @[act.scala 124:19 129:19]
  assign actfunc_io_cfg_act_range_3 = alu_act_param_select_io_cfg_act_range_3; // @[act.scala 124:19 129:19]
  assign actfunc_io_cfg_act_func_prop = alu_act_param_select_io_cfg_act_func_prop; // @[act.scala 124:19 133:23]
  assign actfunc_io_cfg_act_op = io_act_op; // @[act.scala 124:19 125:16]
  assign actfunc_io_cfg_act_en = io_act_en; // @[act.scala 124:19 126:16]
  assign actfunc_io_i_data_data_0 = io_i_data_data_0; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_1 = io_i_data_data_1; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_2 = io_i_data_data_2; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_3 = io_i_data_data_3; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_4 = io_i_data_data_4; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_5 = io_i_data_data_5; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_6 = io_i_data_data_6; // @[act.scala 137:23]
  assign actfunc_io_i_data_data_7 = io_i_data_data_7; // @[act.scala 137:23]
endmodule
module Accel_all(
  input         clock,
  input         reset,
  output        io_resize_load,
  output        io_yolo_finish,
  output        io_conv_finish,
  output [31:0] io_dma_raddr,
  output        io_dma_rareq,
  output [15:0] io_dma_rsize,
  input         io_dma_rbusy,
  input  [63:0] io_dma_rdata,
  input         io_dma_rvalid,
  output        io_dma_rready,
  output [31:0] io_dma_waddr,
  output        io_dma_wareq,
  output [15:0] io_dma_wsize,
  input         io_dma_wbusy,
  output [63:0] io_dma_wdata,
  output        io_dma_wvalid,
  input         io_dma_wready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  control_clock; // @[Accel_all.scala 220:25]
  wire  control_reset; // @[Accel_all.scala 220:25]
  wire  control_io_ap_done; // @[Accel_all.scala 220:25]
  wire  control_io_pool_finish_edge; // @[Accel_all.scala 220:25]
  wire  control_io_conv_finish; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg0; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg1; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg2; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg3; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg4; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg5; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg6; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg7; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg8; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg9; // @[Accel_all.scala 220:25]
  wire [31:0] control_io_reg10; // @[Accel_all.scala 220:25]
  wire  control_io_yolo_finish; // @[Accel_all.scala 220:25]
  wire  control_io_resize_load; // @[Accel_all.scala 220:25]
  wire  control_signal_clock; // @[Accel_all.scala 242:32]
  wire  control_signal_reset; // @[Accel_all.scala 242:32]
  wire  control_signal_io_shutdown; // @[Accel_all.scala 242:32]
  wire  control_signal_io_skip_act; // @[Accel_all.scala 242:32]
  wire [9:0] control_signal_io_conv_col; // @[Accel_all.scala 242:32]
  wire [9:0] control_signal_io_conv_row; // @[Accel_all.scala 242:32]
  wire  control_signal_io_s_mod; // @[Accel_all.scala 242:32]
  wire  control_signal_io_kernal; // @[Accel_all.scala 242:32]
  wire [10:0] control_signal_io_ifmbuf_bram_addr_read_s1; // @[Accel_all.scala 242:32]
  wire  control_signal_io_ifmbuf_addr_read_sel_s1; // @[Accel_all.scala 242:32]
  wire [9:0] control_signal_io_ifmbuf_bram_addr_read_s2_singal; // @[Accel_all.scala 242:32]
  wire [9:0] control_signal_io_ifmbuf_bram_addr_read_s2_double; // @[Accel_all.scala 242:32]
  wire [11:0] control_signal_io_acc_read_addr; // @[Accel_all.scala 242:32]
  wire [11:0] control_signal_io_acc_write_addr; // @[Accel_all.scala 242:32]
  wire  control_signal_io_acc_read_en; // @[Accel_all.scala 242:32]
  wire  control_signal_io_acc_write_en; // @[Accel_all.scala 242:32]
  wire  control_signal_io_acc_curr_data_zero; // @[Accel_all.scala 242:32]
  wire [11:0] control_signal_io_ofm_addr; // @[Accel_all.scala 242:32]
  wire  control_signal_io_ofm_valid; // @[Accel_all.scala 242:32]
  wire  control_signal_io_ofm_done; // @[Accel_all.scala 242:32]
  wire  control_signal_io_pad_top; // @[Accel_all.scala 242:32]
  wire  control_signal_io_pad_bottom; // @[Accel_all.scala 242:32]
  wire  control_signal_io_pad_left_and_right; // @[Accel_all.scala 242:32]
  wire  control_signal_io_pad_size; // @[Accel_all.scala 242:32]
  wire  control_signal_io_zero_pad_valid_s1; // @[Accel_all.scala 242:32]
  wire [4:0] control_signal_io_zero_pad_valid_s2; // @[Accel_all.scala 242:32]
  wire  dma_accel2ddr_clock; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_reset; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_send_enable; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_send_done; // @[Accel_all.scala 271:31]
  wire [31:0] dma_accel2ddr_io_dma_addr; // @[Accel_all.scala 271:31]
  wire [15:0] dma_accel2ddr_io_dma_len; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_dma_wvalid; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_dma_wbusy; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_dma_wready; // @[Accel_all.scala 271:31]
  wire  dma_accel2ddr_io_dma_wareq; // @[Accel_all.scala 271:31]
  wire [31:0] dma_accel2ddr_io_dma_waddr; // @[Accel_all.scala 271:31]
  wire [15:0] dma_accel2ddr_io_dma_wsize; // @[Accel_all.scala 271:31]
  wire [63:0] dma_accel2ddr_io_dma_wdata; // @[Accel_all.scala 271:31]
  wire [16:0] dma_accel2ddr_io_addr_start; // @[Accel_all.scala 271:31]
  wire [16:0] dma_accel2ddr_io_addr_end; // @[Accel_all.scala 271:31]
  wire [16:0] dma_accel2ddr_io_read_addr; // @[Accel_all.scala 271:31]
  wire [63:0] dma_accel2ddr_io_read_data; // @[Accel_all.scala 271:31]
  wire  dma_ddr2accel_clock; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_reset; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_recv_enable; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_recv_done; // @[Accel_all.scala 290:31]
  wire [31:0] dma_ddr2accel_io_dma_addr; // @[Accel_all.scala 290:31]
  wire [15:0] dma_ddr2accel_io_dma_len; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_dma_rvalid; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_dma_rbusy; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_dma_rareq; // @[Accel_all.scala 290:31]
  wire [31:0] dma_ddr2accel_io_dma_raddr; // @[Accel_all.scala 290:31]
  wire [15:0] dma_ddr2accel_io_dma_rsize; // @[Accel_all.scala 290:31]
  wire [63:0] dma_ddr2accel_io_dma_rdata; // @[Accel_all.scala 290:31]
  wire [63:0] dma_ddr2accel_io_write_data; // @[Accel_all.scala 290:31]
  wire  dma_ddr2accel_io_write_enable; // @[Accel_all.scala 290:31]
  wire  generate_ctrl_signal_clock; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_reset; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_recv_enable; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_send_enable; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_conv_start; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_bottleneck_add_enable; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_recv_done; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_send_done; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_conv_done; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_bottleneck_add_done; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_conv_shutdown; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_task_valid; // @[Accel_all.scala 306:38]
  wire  generate_ctrl_signal_io_ap_done; // @[Accel_all.scala 306:38]
  wire [1:0] axis_buf_sel_m_io_axis_buf_sel; // @[Accel_all.scala 322:32]
  wire [63:0] axis_buf_sel_m_io_write_data; // @[Accel_all.scala 322:32]
  wire  axis_buf_sel_m_io_write_enable; // @[Accel_all.scala 322:32]
  wire [63:0] axis_buf_sel_m_io_write_data_ifm; // @[Accel_all.scala 322:32]
  wire  axis_buf_sel_m_io_write_enable_ifm; // @[Accel_all.scala 322:32]
  wire [63:0] axis_buf_sel_m_io_write_data_weight; // @[Accel_all.scala 322:32]
  wire  axis_buf_sel_m_io_write_enable_weight; // @[Accel_all.scala 322:32]
  wire [63:0] axis_buf_sel_m_io_write_data_bias; // @[Accel_all.scala 322:32]
  wire  axis_buf_sel_m_io_write_enable_bias; // @[Accel_all.scala 322:32]
  wire  accel_top_clock; // @[Accel_all.scala 377:27]
  wire  accel_top_reset; // @[Accel_all.scala 377:27]
  wire [2:0] accel_top_io_sel; // @[Accel_all.scala 377:27]
  wire [10:0] accel_top_io_ifmbuf_bram_addr_read_s1; // @[Accel_all.scala 377:27]
  wire  accel_top_io_ifmbuf_bram_addr_read_sel_s1; // @[Accel_all.scala 377:27]
  wire [9:0] accel_top_io_ifmbuf_bram_addr_read_s2_singal; // @[Accel_all.scala 377:27]
  wire [9:0] accel_top_io_ifmbuf_bram_addr_read_s2_double; // @[Accel_all.scala 377:27]
  wire  accel_top_io_ifmbuf_sel; // @[Accel_all.scala 377:27]
  wire  accel_top_io_ifmbuf_bram_en_write; // @[Accel_all.scala 377:27]
  wire  accel_top_io_recv_done; // @[Accel_all.scala 377:27]
  wire  accel_top_io_weightbuf_waddr_clear; // @[Accel_all.scala 377:27]
  wire  accel_top_io_weightbuf_bram_en_write; // @[Accel_all.scala 377:27]
  wire [6:0] accel_top_io_weightbuf_read_addr; // @[Accel_all.scala 377:27]
  wire  accel_top_io_kernal; // @[Accel_all.scala 377:27]
  wire [2:0] accel_top_io_weight_sel; // @[Accel_all.scala 377:27]
  wire  accel_top_io_biasbuf_waddr_clear; // @[Accel_all.scala 377:27]
  wire  accel_top_io_biasbuf_bram_en_write; // @[Accel_all.scala 377:27]
  wire [6:0] accel_top_io_biasbuf_read_addr; // @[Accel_all.scala 377:27]
  wire  accel_top_io_acc_read_en; // @[Accel_all.scala 377:27]
  wire  accel_top_io_acc_write_en; // @[Accel_all.scala 377:27]
  wire [11:0] accel_top_io_acc_read_addr; // @[Accel_all.scala 377:27]
  wire [11:0] accel_top_io_acc_write_addr; // @[Accel_all.scala 377:27]
  wire  accel_top_io_acc_prev_data_zero; // @[Accel_all.scala 377:27]
  wire  accel_top_io_acc_curr_data_zero; // @[Accel_all.scala 377:27]
  wire  accel_top_io_ofmbuf_bram_en_write; // @[Accel_all.scala 377:27]
  wire [11:0] accel_top_io_ofmbuf_bram_write_addr; // @[Accel_all.scala 377:27]
  wire [63:0] accel_top_io_ofmbuf_bram_read_addr; // @[Accel_all.scala 377:27]
  wire [9:0] accel_top_io_col; // @[Accel_all.scala 377:27]
  wire [9:0] accel_top_io_row; // @[Accel_all.scala 377:27]
  wire  accel_top_io_pad_top; // @[Accel_all.scala 377:27]
  wire  accel_top_io_pad_bottom; // @[Accel_all.scala 377:27]
  wire  accel_top_io_pad_left_and_right; // @[Accel_all.scala 377:27]
  wire [4:0] accel_top_io_zero_pad_valid_s2; // @[Accel_all.scala 377:27]
  wire  accel_top_io_zero_pad_valid_s1; // @[Accel_all.scala 377:27]
  wire [15:0] accel_top_io_scale; // @[Accel_all.scala 377:27]
  wire [3:0] accel_top_io_shift; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_zero_point_in; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_zero_point_out; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_zero_point_A_act; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_ifm_in_7; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_weight_in_7; // @[Accel_all.scala 377:27]
  wire [17:0] accel_top_io_bias_in; // @[Accel_all.scala 377:27]
  wire  accel_top_io_bias_valid; // @[Accel_all.scala 377:27]
  wire [63:0] accel_top_io_ofm_out_bundle; // @[Accel_all.scala 377:27]
  wire  accel_top_io_skip_act; // @[Accel_all.scala 377:27]
  wire  accel_top_io_pool_enable; // @[Accel_all.scala 377:27]
  wire  accel_top_io_pool_finish; // @[Accel_all.scala 377:27]
  wire  accel_top_io_upsample_enable; // @[Accel_all.scala 377:27]
  wire  accel_top_io_bottleneck_add_enable; // @[Accel_all.scala 377:27]
  wire  accel_top_io_bottleneck_add_finish; // @[Accel_all.scala 377:27]
  wire  accel_top_io_s_mod; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_indata_7; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_act_outdata_7; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in0_7; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_in1_7; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_0; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_1; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_2; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_3; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_4; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_5; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_6; // @[Accel_all.scala 377:27]
  wire [7:0] accel_top_io_bn_add_result_7; // @[Accel_all.scala 377:27]
  wire  accel_top_io_yolo_cls_en; // @[Accel_all.scala 377:27]
  wire [63:0] accel_top_io_yolo_cls_data_before_compare; // @[Accel_all.scala 377:27]
  wire [63:0] accel_top_io_yolo_cls_data_after_compare; // @[Accel_all.scala 377:27]
  wire  yolo_clock; // @[Accel_all.scala 464:22]
  wire  yolo_reset; // @[Accel_all.scala 464:22]
  wire  yolo_io_yolo_layer_cls_en; // @[Accel_all.scala 464:22]
  wire  yolo_io_yolo_cls_finish; // @[Accel_all.scala 464:22]
  wire [1:0] yolo_io_yolo_current_cls_detect_layer; // @[Accel_all.scala 464:22]
  wire [3:0] yolo_io_yolo_layer_cls_div_cnt; // @[Accel_all.scala 464:22]
  wire [11:0] yolo_io_ofm_read_addr; // @[Accel_all.scala 464:22]
  wire [63:0] yolo_io_ofm_write_data_before; // @[Accel_all.scala 464:22]
  wire  yolo_io_ofm_write_en_before; // @[Accel_all.scala 464:22]
  wire [63:0] yolo_io_ofm_write_data_after; // @[Accel_all.scala 464:22]
  wire  yolo_io_ofm_write_en_after; // @[Accel_all.scala 464:22]
  wire [11:0] yolo_io_ofm_write_addr_after; // @[Accel_all.scala 464:22]
  wire [7:0] yolo_io_data_before_sigmoid; // @[Accel_all.scala 464:22]
  wire [23:0] yolo_io_data_after_sigmoid; // @[Accel_all.scala 464:22]
  wire  yolo_io_sigmoid_en; // @[Accel_all.scala 464:22]
  wire  dequant_clock; // @[Accel_all.scala 494:25]
  wire  dequant_reset; // @[Accel_all.scala 494:25]
  wire  dequant_io_en; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_0; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_1; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_2; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_3; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_4; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_5; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_6; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_i_data_7; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_scale; // @[Accel_all.scala 494:25]
  wire [7:0] dequant_io_zero_point; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_0; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_1; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_2; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_3; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_4; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_5; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_6; // @[Accel_all.scala 494:25]
  wire [31:0] dequant_io_o_data_7; // @[Accel_all.scala 494:25]
  wire  dequant_extra_clock; // @[Accel_all.scala 501:31]
  wire  dequant_extra_reset; // @[Accel_all.scala 501:31]
  wire  dequant_extra_io_en; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_0; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_1; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_2; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_3; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_4; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_5; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_6; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_i_data_7; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_scale; // @[Accel_all.scala 501:31]
  wire [7:0] dequant_extra_io_zero_point; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_0; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_1; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_2; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_3; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_4; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_5; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_6; // @[Accel_all.scala 501:31]
  wire [31:0] dequant_extra_io_o_data_7; // @[Accel_all.scala 501:31]
  wire  bn_add_float_result_0_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_0_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_0_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_0_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_0_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_0_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_1_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_1_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_1_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_1_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_1_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_1_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_2_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_2_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_2_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_2_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_2_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_2_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_3_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_3_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_3_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_3_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_3_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_3_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_4_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_4_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_4_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_4_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_4_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_4_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_5_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_5_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_5_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_5_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_5_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_5_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_6_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_6_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_6_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_6_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_6_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_6_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_7_adder_clock; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_7_adder_reset; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_7_adder_io_x; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_7_adder_io_y; // @[Arithmetic.scala 115:25]
  wire [31:0] bn_add_float_result_7_adder_io_z; // @[Arithmetic.scala 115:25]
  wire  bn_add_float_result_7_adder_io_valid_in; // @[Arithmetic.scala 115:25]
  wire  quant_clock; // @[Accel_all.scala 514:23]
  wire  quant_reset; // @[Accel_all.scala 514:23]
  wire  quant_io_en; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_0; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_1; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_2; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_3; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_4; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_5; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_6; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_i_data_7; // @[Accel_all.scala 514:23]
  wire [31:0] quant_io_scale; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_zero_point; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_0; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_1; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_2; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_3; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_4; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_5; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_6; // @[Accel_all.scala 514:23]
  wire [7:0] quant_io_o_data_7; // @[Accel_all.scala 514:23]
  wire  alu_act_clock; // @[Accel_all.scala 522:25]
  wire  alu_act_reset; // @[Accel_all.scala 522:25]
  wire [1:0] alu_act_io_act_op; // @[Accel_all.scala 522:25]
  wire  alu_act_io_act_en; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_0; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_1; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_2; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_3; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_4; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_5; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_6; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_i_data_data_7; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_0; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_1; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_2; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_3; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_4; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_5; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_6; // @[Accel_all.scala 522:25]
  wire [31:0] alu_act_io_o_data_data_7; // @[Accel_all.scala 522:25]
  wire [31:0] reg_8 = control_io_reg8; // @[Accel_all.scala 232:10 53:21]
  wire  yolo_cls_en = reg_8[16]; // @[Accel_all.scala 179:25]
  wire  yolo_cls_finish = yolo_io_yolo_cls_finish; // @[Accel_all.scala 466:21 98:31]
  wire  ofm_done = control_signal_io_ofm_done; // @[Accel_all.scala 113:24 261:13]
  wire [31:0] reg_0 = control_io_reg0; // @[Accel_all.scala 224:10 43:21]
  wire  pool_enable = reg_0[5]; // @[Accel_all.scala 132:25]
  wire  task_valid = reg_0[9]; // @[Accel_all.scala 136:24]
  wire [2:0] pad_cfg = reg_0[15:13]; // @[Accel_all.scala 138:21]
  wire  skip_act = reg_0[17]; // @[Accel_all.scala 140:20]
  wire [7:0] row = reg_0[31:24]; // @[Accel_all.scala 144:20]
  wire [31:0] reg_1 = control_io_reg1; // @[Accel_all.scala 225:10 44:21]
  wire [31:0] reg_2 = control_io_reg2; // @[Accel_all.scala 226:10 45:21]
  wire [7:0] dequant_zero_point = reg_2[15:8]; // @[Accel_all.scala 151:31]
  reg  weightbuf_waddr_clear_REG; // @[utils.scala 10:17]
  reg  biasbuf_waddr_clear_REG; // @[utils.scala 10:17]
  wire [31:0] reg_3 = control_io_reg3; // @[Accel_all.scala 227:10 46:21]
  wire [31:0] reg_5 = control_io_reg5; // @[Accel_all.scala 229:10 49:21]
  wire [31:0] reg_7 = control_io_reg7; // @[Accel_all.scala 231:10 51:21]
  wire [15:0] dma_accel2ddr_len = reg_7[18:3]; // @[Accel_all.scala 170:35]
  wire [1:0] pool_cnt = reg_8[11:10]; // @[Accel_all.scala 178:22]
  wire  ofm_write_disable = reg_8[17]; // @[Accel_all.scala 180:31]
  reg [31:0] dequant_extra_scala_temp; // @[Reg.scala 35:20]
  wire  conv_finish_from_control = control_io_conv_finish; // @[Accel_all.scala 189:40 223:29]
  wire [31:0] dequant_scala = control_io_reg9; // @[Accel_all.scala 233:10 54:21]
  reg [31:0] dequant_extra_scala; // @[Reg.scala 35:20]
  reg [7:0] dequant_extra_zero_point_temp; // @[Reg.scala 35:20]
  reg [7:0] dequant_extra_zero_point; // @[Reg.scala 35:20]
  wire [10:0] _addr_start_T = pool_cnt * 9'h190; // @[Accel_all.scala 199:45]
  wire [10:0] _addr_start_T_1 = pool_enable ? _addr_start_T : 11'h0; // @[Accel_all.scala 199:22]
  wire [15:0] addr_start = {{5'd0}, _addr_start_T_1}; // @[Accel_all.scala 199:16 62:26]
  wire [15:0] addr_end = dma_accel2ddr_len + addr_start; // @[Accel_all.scala 200:35]
  wire [63:0] write_data_ifm = axis_buf_sel_m_io_write_data_ifm; // @[Accel_all.scala 328:20 79:30]
  wire [63:0] write_data_weight = axis_buf_sel_m_io_write_data_weight; // @[Accel_all.scala 331:23 82:33]
  wire [15:0] read_addr = dma_accel2ddr_io_read_addr[15:0]; // @[Accel_all.scala 288:15 64:25]
  wire [11:0] ofmbuf_bram_read_addr = read_addr[11:0]; // @[Accel_all.scala 353:37]
  wire  yolo_ofm_write_en_after = yolo_io_ofm_write_en_after; // @[Accel_all.scala 368:37 475:29]
  wire  ofm_valid = control_signal_io_ofm_valid; // @[Accel_all.scala 112:25 260:14]
  wire [63:0] yolo_ofm_write_addr_after = {{52'd0}, yolo_io_ofm_write_addr_after}; // @[Accel_all.scala 369:39 476:31]
  wire [11:0] ofm_addr = control_signal_io_ofm_addr; // @[Accel_all.scala 111:24 259:13]
  wire [63:0] _accel_top_io_ofmbuf_bram_write_addr_T = yolo_cls_en ? yolo_ofm_write_addr_after : {{52'd0}, ofm_addr}; // @[Accel_all.scala 409:47]
  wire [11:0] yolo_ofm_read_addr = yolo_io_ofm_read_addr; // @[Accel_all.scala 366:32 470:24]
  wire [11:0] _accel_top_io_ofmbuf_bram_read_addr_T = yolo_cls_en ? yolo_ofm_read_addr : ofmbuf_bram_read_addr; // @[Accel_all.scala 410:46]
  wire  _act_op_T = ~skip_act; // @[Accel_all.scala 463:41]
  wire  sigmoid_en = yolo_io_sigmoid_en; // @[Accel_all.scala 462:24 477:15]
  wire [31:0] alu_act_out_0 = alu_act_io_o_data_data_0; // @[Accel_all.scala 375:27 525:17]
  wire  bn_add_working = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  wire [7:0] yolo_data_before_sigmoid = yolo_io_data_before_sigmoid; // @[Accel_all.scala 372:40 478:30]
  wire [7:0] _dequant_in_0_T_3 = sigmoid_en ? yolo_data_before_sigmoid : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] bn_add_in0_0 = accel_top_io_bn_add_in0_0; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_0_T_4 = bn_add_working ? bn_add_in0_0 : _dequant_in_0_T_3; // @[Mux.scala 101:16]
  wire [7:0] act_indata_0 = accel_top_io_act_indata_0; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_1 = accel_top_io_bn_add_in0_1; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_1_T_2 = bn_add_working ? bn_add_in0_1 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_1 = accel_top_io_act_indata_1; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_2 = accel_top_io_bn_add_in0_2; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_2_T_2 = bn_add_working ? bn_add_in0_2 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_2 = accel_top_io_act_indata_2; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_3 = accel_top_io_bn_add_in0_3; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_3_T_2 = bn_add_working ? bn_add_in0_3 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_3 = accel_top_io_act_indata_3; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_4 = accel_top_io_bn_add_in0_4; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_4_T_2 = bn_add_working ? bn_add_in0_4 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_4 = accel_top_io_act_indata_4; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_5 = accel_top_io_bn_add_in0_5; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_5_T_2 = bn_add_working ? bn_add_in0_5 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_5 = accel_top_io_act_indata_5; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_6 = accel_top_io_bn_add_in0_6; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_6_T_2 = bn_add_working ? bn_add_in0_6 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_6 = accel_top_io_act_indata_6; // @[Accel_all.scala 356:26 421:20]
  wire [7:0] bn_add_in0_7 = accel_top_io_bn_add_in0_7; // @[Accel_all.scala 358:26 452:16]
  wire [7:0] _dequant_in_7_T_2 = bn_add_working ? bn_add_in0_7 : 8'h0; // @[Mux.scala 101:16]
  wire [7:0] act_indata_7 = accel_top_io_act_indata_7; // @[Accel_all.scala 356:26 421:20]
  wire [31:0] bn_add_float_result_0_result_2_bits = bn_add_float_result_0_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] bn_add_float_result_1_result_2_bits = bn_add_float_result_1_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_1 = alu_act_io_o_data_data_1; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_2_result_2_bits = bn_add_float_result_2_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_2 = alu_act_io_o_data_data_2; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_3_result_2_bits = bn_add_float_result_3_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_3 = alu_act_io_o_data_data_3; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_4_result_2_bits = bn_add_float_result_4_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_4 = alu_act_io_o_data_data_4; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_5_result_2_bits = bn_add_float_result_5_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_5 = alu_act_io_o_data_data_5; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_6_result_2_bits = bn_add_float_result_6_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_6 = alu_act_io_o_data_data_6; // @[Accel_all.scala 375:27 525:17]
  wire [31:0] bn_add_float_result_7_result_2_bits = bn_add_float_result_7_adder_io_z; // @[Arithmetic.scala 124:22 125:17]
  wire [31:0] alu_act_out_7 = alu_act_io_o_data_data_7; // @[Accel_all.scala 375:27 525:17]
  wire [63:0] write_data_bias = axis_buf_sel_m_io_write_data_bias; // @[Accel_all.scala 334:21 85:31]
  accel_control control ( // @[Accel_all.scala 220:25]
    .clock(control_clock),
    .reset(control_reset),
    .io_ap_done(control_io_ap_done),
    .io_pool_finish_edge(control_io_pool_finish_edge),
    .io_conv_finish(control_io_conv_finish),
    .io_reg0(control_io_reg0),
    .io_reg1(control_io_reg1),
    .io_reg2(control_io_reg2),
    .io_reg3(control_io_reg3),
    .io_reg4(control_io_reg4),
    .io_reg5(control_io_reg5),
    .io_reg6(control_io_reg6),
    .io_reg7(control_io_reg7),
    .io_reg8(control_io_reg8),
    .io_reg9(control_io_reg9),
    .io_reg10(control_io_reg10),
    .io_yolo_finish(control_io_yolo_finish),
    .io_resize_load(control_io_resize_load)
  );
  control_signal control_signal ( // @[Accel_all.scala 242:32]
    .clock(control_signal_clock),
    .reset(control_signal_reset),
    .io_shutdown(control_signal_io_shutdown),
    .io_skip_act(control_signal_io_skip_act),
    .io_conv_col(control_signal_io_conv_col),
    .io_conv_row(control_signal_io_conv_row),
    .io_s_mod(control_signal_io_s_mod),
    .io_kernal(control_signal_io_kernal),
    .io_ifmbuf_bram_addr_read_s1(control_signal_io_ifmbuf_bram_addr_read_s1),
    .io_ifmbuf_addr_read_sel_s1(control_signal_io_ifmbuf_addr_read_sel_s1),
    .io_ifmbuf_bram_addr_read_s2_singal(control_signal_io_ifmbuf_bram_addr_read_s2_singal),
    .io_ifmbuf_bram_addr_read_s2_double(control_signal_io_ifmbuf_bram_addr_read_s2_double),
    .io_acc_read_addr(control_signal_io_acc_read_addr),
    .io_acc_write_addr(control_signal_io_acc_write_addr),
    .io_acc_read_en(control_signal_io_acc_read_en),
    .io_acc_write_en(control_signal_io_acc_write_en),
    .io_acc_curr_data_zero(control_signal_io_acc_curr_data_zero),
    .io_ofm_addr(control_signal_io_ofm_addr),
    .io_ofm_valid(control_signal_io_ofm_valid),
    .io_ofm_done(control_signal_io_ofm_done),
    .io_pad_top(control_signal_io_pad_top),
    .io_pad_bottom(control_signal_io_pad_bottom),
    .io_pad_left_and_right(control_signal_io_pad_left_and_right),
    .io_pad_size(control_signal_io_pad_size),
    .io_zero_pad_valid_s1(control_signal_io_zero_pad_valid_s1),
    .io_zero_pad_valid_s2(control_signal_io_zero_pad_valid_s2)
  );
  DMA_Master dma_accel2ddr ( // @[Accel_all.scala 271:31]
    .clock(dma_accel2ddr_clock),
    .reset(dma_accel2ddr_reset),
    .io_send_enable(dma_accel2ddr_io_send_enable),
    .io_send_done(dma_accel2ddr_io_send_done),
    .io_dma_addr(dma_accel2ddr_io_dma_addr),
    .io_dma_len(dma_accel2ddr_io_dma_len),
    .io_dma_wvalid(dma_accel2ddr_io_dma_wvalid),
    .io_dma_wbusy(dma_accel2ddr_io_dma_wbusy),
    .io_dma_wready(dma_accel2ddr_io_dma_wready),
    .io_dma_wareq(dma_accel2ddr_io_dma_wareq),
    .io_dma_waddr(dma_accel2ddr_io_dma_waddr),
    .io_dma_wsize(dma_accel2ddr_io_dma_wsize),
    .io_dma_wdata(dma_accel2ddr_io_dma_wdata),
    .io_addr_start(dma_accel2ddr_io_addr_start),
    .io_addr_end(dma_accel2ddr_io_addr_end),
    .io_read_addr(dma_accel2ddr_io_read_addr),
    .io_read_data(dma_accel2ddr_io_read_data)
  );
  DMA_Slave dma_ddr2accel ( // @[Accel_all.scala 290:31]
    .clock(dma_ddr2accel_clock),
    .reset(dma_ddr2accel_reset),
    .io_recv_enable(dma_ddr2accel_io_recv_enable),
    .io_recv_done(dma_ddr2accel_io_recv_done),
    .io_dma_addr(dma_ddr2accel_io_dma_addr),
    .io_dma_len(dma_ddr2accel_io_dma_len),
    .io_dma_rvalid(dma_ddr2accel_io_dma_rvalid),
    .io_dma_rbusy(dma_ddr2accel_io_dma_rbusy),
    .io_dma_rareq(dma_ddr2accel_io_dma_rareq),
    .io_dma_raddr(dma_ddr2accel_io_dma_raddr),
    .io_dma_rsize(dma_ddr2accel_io_dma_rsize),
    .io_dma_rdata(dma_ddr2accel_io_dma_rdata),
    .io_write_data(dma_ddr2accel_io_write_data),
    .io_write_enable(dma_ddr2accel_io_write_enable)
  );
  generate_ctrl_signal generate_ctrl_signal ( // @[Accel_all.scala 306:38]
    .clock(generate_ctrl_signal_clock),
    .reset(generate_ctrl_signal_reset),
    .io_recv_enable(generate_ctrl_signal_io_recv_enable),
    .io_send_enable(generate_ctrl_signal_io_send_enable),
    .io_conv_start(generate_ctrl_signal_io_conv_start),
    .io_bottleneck_add_enable(generate_ctrl_signal_io_bottleneck_add_enable),
    .io_recv_done(generate_ctrl_signal_io_recv_done),
    .io_send_done(generate_ctrl_signal_io_send_done),
    .io_conv_done(generate_ctrl_signal_io_conv_done),
    .io_bottleneck_add_done(generate_ctrl_signal_io_bottleneck_add_done),
    .io_conv_shutdown(generate_ctrl_signal_io_conv_shutdown),
    .io_bn_add_working(generate_ctrl_signal_io_bn_add_working),
    .io_task_valid(generate_ctrl_signal_io_task_valid),
    .io_ap_done(generate_ctrl_signal_io_ap_done)
  );
  axis_buf_sel axis_buf_sel_m ( // @[Accel_all.scala 322:32]
    .io_axis_buf_sel(axis_buf_sel_m_io_axis_buf_sel),
    .io_write_data(axis_buf_sel_m_io_write_data),
    .io_write_enable(axis_buf_sel_m_io_write_enable),
    .io_write_data_ifm(axis_buf_sel_m_io_write_data_ifm),
    .io_write_enable_ifm(axis_buf_sel_m_io_write_enable_ifm),
    .io_write_data_weight(axis_buf_sel_m_io_write_data_weight),
    .io_write_enable_weight(axis_buf_sel_m_io_write_enable_weight),
    .io_write_data_bias(axis_buf_sel_m_io_write_data_bias),
    .io_write_enable_bias(axis_buf_sel_m_io_write_enable_bias)
  );
  accel_top accel_top ( // @[Accel_all.scala 377:27]
    .clock(accel_top_clock),
    .reset(accel_top_reset),
    .io_sel(accel_top_io_sel),
    .io_ifmbuf_bram_addr_read_s1(accel_top_io_ifmbuf_bram_addr_read_s1),
    .io_ifmbuf_bram_addr_read_sel_s1(accel_top_io_ifmbuf_bram_addr_read_sel_s1),
    .io_ifmbuf_bram_addr_read_s2_singal(accel_top_io_ifmbuf_bram_addr_read_s2_singal),
    .io_ifmbuf_bram_addr_read_s2_double(accel_top_io_ifmbuf_bram_addr_read_s2_double),
    .io_ifmbuf_sel(accel_top_io_ifmbuf_sel),
    .io_ifmbuf_bram_en_write(accel_top_io_ifmbuf_bram_en_write),
    .io_recv_done(accel_top_io_recv_done),
    .io_weightbuf_waddr_clear(accel_top_io_weightbuf_waddr_clear),
    .io_weightbuf_bram_en_write(accel_top_io_weightbuf_bram_en_write),
    .io_weightbuf_read_addr(accel_top_io_weightbuf_read_addr),
    .io_kernal(accel_top_io_kernal),
    .io_weight_sel(accel_top_io_weight_sel),
    .io_biasbuf_waddr_clear(accel_top_io_biasbuf_waddr_clear),
    .io_biasbuf_bram_en_write(accel_top_io_biasbuf_bram_en_write),
    .io_biasbuf_read_addr(accel_top_io_biasbuf_read_addr),
    .io_acc_read_en(accel_top_io_acc_read_en),
    .io_acc_write_en(accel_top_io_acc_write_en),
    .io_acc_read_addr(accel_top_io_acc_read_addr),
    .io_acc_write_addr(accel_top_io_acc_write_addr),
    .io_acc_prev_data_zero(accel_top_io_acc_prev_data_zero),
    .io_acc_curr_data_zero(accel_top_io_acc_curr_data_zero),
    .io_ofmbuf_bram_en_write(accel_top_io_ofmbuf_bram_en_write),
    .io_ofmbuf_bram_write_addr(accel_top_io_ofmbuf_bram_write_addr),
    .io_ofmbuf_bram_read_addr(accel_top_io_ofmbuf_bram_read_addr),
    .io_col(accel_top_io_col),
    .io_row(accel_top_io_row),
    .io_pad_top(accel_top_io_pad_top),
    .io_pad_bottom(accel_top_io_pad_bottom),
    .io_pad_left_and_right(accel_top_io_pad_left_and_right),
    .io_zero_pad_valid_s2(accel_top_io_zero_pad_valid_s2),
    .io_zero_pad_valid_s1(accel_top_io_zero_pad_valid_s1),
    .io_scale(accel_top_io_scale),
    .io_shift(accel_top_io_shift),
    .io_zero_point_in(accel_top_io_zero_point_in),
    .io_zero_point_out(accel_top_io_zero_point_out),
    .io_zero_point_A_act(accel_top_io_zero_point_A_act),
    .io_ifm_in_0(accel_top_io_ifm_in_0),
    .io_ifm_in_1(accel_top_io_ifm_in_1),
    .io_ifm_in_2(accel_top_io_ifm_in_2),
    .io_ifm_in_3(accel_top_io_ifm_in_3),
    .io_ifm_in_4(accel_top_io_ifm_in_4),
    .io_ifm_in_5(accel_top_io_ifm_in_5),
    .io_ifm_in_6(accel_top_io_ifm_in_6),
    .io_ifm_in_7(accel_top_io_ifm_in_7),
    .io_weight_in_0(accel_top_io_weight_in_0),
    .io_weight_in_1(accel_top_io_weight_in_1),
    .io_weight_in_2(accel_top_io_weight_in_2),
    .io_weight_in_3(accel_top_io_weight_in_3),
    .io_weight_in_4(accel_top_io_weight_in_4),
    .io_weight_in_5(accel_top_io_weight_in_5),
    .io_weight_in_6(accel_top_io_weight_in_6),
    .io_weight_in_7(accel_top_io_weight_in_7),
    .io_bias_in(accel_top_io_bias_in),
    .io_bias_valid(accel_top_io_bias_valid),
    .io_ofm_out_bundle(accel_top_io_ofm_out_bundle),
    .io_skip_act(accel_top_io_skip_act),
    .io_pool_enable(accel_top_io_pool_enable),
    .io_pool_finish(accel_top_io_pool_finish),
    .io_upsample_enable(accel_top_io_upsample_enable),
    .io_bottleneck_add_enable(accel_top_io_bottleneck_add_enable),
    .io_bottleneck_add_finish(accel_top_io_bottleneck_add_finish),
    .io_s_mod(accel_top_io_s_mod),
    .io_act_indata_0(accel_top_io_act_indata_0),
    .io_act_indata_1(accel_top_io_act_indata_1),
    .io_act_indata_2(accel_top_io_act_indata_2),
    .io_act_indata_3(accel_top_io_act_indata_3),
    .io_act_indata_4(accel_top_io_act_indata_4),
    .io_act_indata_5(accel_top_io_act_indata_5),
    .io_act_indata_6(accel_top_io_act_indata_6),
    .io_act_indata_7(accel_top_io_act_indata_7),
    .io_act_outdata_0(accel_top_io_act_outdata_0),
    .io_act_outdata_1(accel_top_io_act_outdata_1),
    .io_act_outdata_2(accel_top_io_act_outdata_2),
    .io_act_outdata_3(accel_top_io_act_outdata_3),
    .io_act_outdata_4(accel_top_io_act_outdata_4),
    .io_act_outdata_5(accel_top_io_act_outdata_5),
    .io_act_outdata_6(accel_top_io_act_outdata_6),
    .io_act_outdata_7(accel_top_io_act_outdata_7),
    .io_bn_add_in0_0(accel_top_io_bn_add_in0_0),
    .io_bn_add_in0_1(accel_top_io_bn_add_in0_1),
    .io_bn_add_in0_2(accel_top_io_bn_add_in0_2),
    .io_bn_add_in0_3(accel_top_io_bn_add_in0_3),
    .io_bn_add_in0_4(accel_top_io_bn_add_in0_4),
    .io_bn_add_in0_5(accel_top_io_bn_add_in0_5),
    .io_bn_add_in0_6(accel_top_io_bn_add_in0_6),
    .io_bn_add_in0_7(accel_top_io_bn_add_in0_7),
    .io_bn_add_in1_0(accel_top_io_bn_add_in1_0),
    .io_bn_add_in1_1(accel_top_io_bn_add_in1_1),
    .io_bn_add_in1_2(accel_top_io_bn_add_in1_2),
    .io_bn_add_in1_3(accel_top_io_bn_add_in1_3),
    .io_bn_add_in1_4(accel_top_io_bn_add_in1_4),
    .io_bn_add_in1_5(accel_top_io_bn_add_in1_5),
    .io_bn_add_in1_6(accel_top_io_bn_add_in1_6),
    .io_bn_add_in1_7(accel_top_io_bn_add_in1_7),
    .io_bn_add_result_0(accel_top_io_bn_add_result_0),
    .io_bn_add_result_1(accel_top_io_bn_add_result_1),
    .io_bn_add_result_2(accel_top_io_bn_add_result_2),
    .io_bn_add_result_3(accel_top_io_bn_add_result_3),
    .io_bn_add_result_4(accel_top_io_bn_add_result_4),
    .io_bn_add_result_5(accel_top_io_bn_add_result_5),
    .io_bn_add_result_6(accel_top_io_bn_add_result_6),
    .io_bn_add_result_7(accel_top_io_bn_add_result_7),
    .io_yolo_cls_en(accel_top_io_yolo_cls_en),
    .io_yolo_cls_data_before_compare(accel_top_io_yolo_cls_data_before_compare),
    .io_yolo_cls_data_after_compare(accel_top_io_yolo_cls_data_after_compare)
  );
  yolo_layer yolo ( // @[Accel_all.scala 464:22]
    .clock(yolo_clock),
    .reset(yolo_reset),
    .io_yolo_layer_cls_en(yolo_io_yolo_layer_cls_en),
    .io_yolo_cls_finish(yolo_io_yolo_cls_finish),
    .io_yolo_current_cls_detect_layer(yolo_io_yolo_current_cls_detect_layer),
    .io_yolo_layer_cls_div_cnt(yolo_io_yolo_layer_cls_div_cnt),
    .io_ofm_read_addr(yolo_io_ofm_read_addr),
    .io_ofm_write_data_before(yolo_io_ofm_write_data_before),
    .io_ofm_write_en_before(yolo_io_ofm_write_en_before),
    .io_ofm_write_data_after(yolo_io_ofm_write_data_after),
    .io_ofm_write_en_after(yolo_io_ofm_write_en_after),
    .io_ofm_write_addr_after(yolo_io_ofm_write_addr_after),
    .io_data_before_sigmoid(yolo_io_data_before_sigmoid),
    .io_data_after_sigmoid(yolo_io_data_after_sigmoid),
    .io_sigmoid_en(yolo_io_sigmoid_en)
  );
  dequant_int8_2_fp32 dequant ( // @[Accel_all.scala 494:25]
    .clock(dequant_clock),
    .reset(dequant_reset),
    .io_en(dequant_io_en),
    .io_i_data_0(dequant_io_i_data_0),
    .io_i_data_1(dequant_io_i_data_1),
    .io_i_data_2(dequant_io_i_data_2),
    .io_i_data_3(dequant_io_i_data_3),
    .io_i_data_4(dequant_io_i_data_4),
    .io_i_data_5(dequant_io_i_data_5),
    .io_i_data_6(dequant_io_i_data_6),
    .io_i_data_7(dequant_io_i_data_7),
    .io_scale(dequant_io_scale),
    .io_zero_point(dequant_io_zero_point),
    .io_o_data_0(dequant_io_o_data_0),
    .io_o_data_1(dequant_io_o_data_1),
    .io_o_data_2(dequant_io_o_data_2),
    .io_o_data_3(dequant_io_o_data_3),
    .io_o_data_4(dequant_io_o_data_4),
    .io_o_data_5(dequant_io_o_data_5),
    .io_o_data_6(dequant_io_o_data_6),
    .io_o_data_7(dequant_io_o_data_7)
  );
  dequant_int8_2_fp32 dequant_extra ( // @[Accel_all.scala 501:31]
    .clock(dequant_extra_clock),
    .reset(dequant_extra_reset),
    .io_en(dequant_extra_io_en),
    .io_i_data_0(dequant_extra_io_i_data_0),
    .io_i_data_1(dequant_extra_io_i_data_1),
    .io_i_data_2(dequant_extra_io_i_data_2),
    .io_i_data_3(dequant_extra_io_i_data_3),
    .io_i_data_4(dequant_extra_io_i_data_4),
    .io_i_data_5(dequant_extra_io_i_data_5),
    .io_i_data_6(dequant_extra_io_i_data_6),
    .io_i_data_7(dequant_extra_io_i_data_7),
    .io_scale(dequant_extra_io_scale),
    .io_zero_point(dequant_extra_io_zero_point),
    .io_o_data_0(dequant_extra_io_o_data_0),
    .io_o_data_1(dequant_extra_io_o_data_1),
    .io_o_data_2(dequant_extra_io_o_data_2),
    .io_o_data_3(dequant_extra_io_o_data_3),
    .io_o_data_4(dequant_extra_io_o_data_4),
    .io_o_data_5(dequant_extra_io_o_data_5),
    .io_o_data_6(dequant_extra_io_o_data_6),
    .io_o_data_7(dequant_extra_io_o_data_7)
  );
  FP32_Adder bn_add_float_result_0_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_0_adder_clock),
    .reset(bn_add_float_result_0_adder_reset),
    .io_x(bn_add_float_result_0_adder_io_x),
    .io_y(bn_add_float_result_0_adder_io_y),
    .io_z(bn_add_float_result_0_adder_io_z),
    .io_valid_in(bn_add_float_result_0_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_1_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_1_adder_clock),
    .reset(bn_add_float_result_1_adder_reset),
    .io_x(bn_add_float_result_1_adder_io_x),
    .io_y(bn_add_float_result_1_adder_io_y),
    .io_z(bn_add_float_result_1_adder_io_z),
    .io_valid_in(bn_add_float_result_1_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_2_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_2_adder_clock),
    .reset(bn_add_float_result_2_adder_reset),
    .io_x(bn_add_float_result_2_adder_io_x),
    .io_y(bn_add_float_result_2_adder_io_y),
    .io_z(bn_add_float_result_2_adder_io_z),
    .io_valid_in(bn_add_float_result_2_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_3_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_3_adder_clock),
    .reset(bn_add_float_result_3_adder_reset),
    .io_x(bn_add_float_result_3_adder_io_x),
    .io_y(bn_add_float_result_3_adder_io_y),
    .io_z(bn_add_float_result_3_adder_io_z),
    .io_valid_in(bn_add_float_result_3_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_4_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_4_adder_clock),
    .reset(bn_add_float_result_4_adder_reset),
    .io_x(bn_add_float_result_4_adder_io_x),
    .io_y(bn_add_float_result_4_adder_io_y),
    .io_z(bn_add_float_result_4_adder_io_z),
    .io_valid_in(bn_add_float_result_4_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_5_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_5_adder_clock),
    .reset(bn_add_float_result_5_adder_reset),
    .io_x(bn_add_float_result_5_adder_io_x),
    .io_y(bn_add_float_result_5_adder_io_y),
    .io_z(bn_add_float_result_5_adder_io_z),
    .io_valid_in(bn_add_float_result_5_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_6_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_6_adder_clock),
    .reset(bn_add_float_result_6_adder_reset),
    .io_x(bn_add_float_result_6_adder_io_x),
    .io_y(bn_add_float_result_6_adder_io_y),
    .io_z(bn_add_float_result_6_adder_io_z),
    .io_valid_in(bn_add_float_result_6_adder_io_valid_in)
  );
  FP32_Adder bn_add_float_result_7_adder ( // @[Arithmetic.scala 115:25]
    .clock(bn_add_float_result_7_adder_clock),
    .reset(bn_add_float_result_7_adder_reset),
    .io_x(bn_add_float_result_7_adder_io_x),
    .io_y(bn_add_float_result_7_adder_io_y),
    .io_z(bn_add_float_result_7_adder_io_z),
    .io_valid_in(bn_add_float_result_7_adder_io_valid_in)
  );
  quant_fp32_2_int8 quant ( // @[Accel_all.scala 514:23]
    .clock(quant_clock),
    .reset(quant_reset),
    .io_en(quant_io_en),
    .io_i_data_0(quant_io_i_data_0),
    .io_i_data_1(quant_io_i_data_1),
    .io_i_data_2(quant_io_i_data_2),
    .io_i_data_3(quant_io_i_data_3),
    .io_i_data_4(quant_io_i_data_4),
    .io_i_data_5(quant_io_i_data_5),
    .io_i_data_6(quant_io_i_data_6),
    .io_i_data_7(quant_io_i_data_7),
    .io_scale(quant_io_scale),
    .io_zero_point(quant_io_zero_point),
    .io_o_data_0(quant_io_o_data_0),
    .io_o_data_1(quant_io_o_data_1),
    .io_o_data_2(quant_io_o_data_2),
    .io_o_data_3(quant_io_o_data_3),
    .io_o_data_4(quant_io_o_data_4),
    .io_o_data_5(quant_io_o_data_5),
    .io_o_data_6(quant_io_o_data_6),
    .io_o_data_7(quant_io_o_data_7)
  );
  alu_act alu_act ( // @[Accel_all.scala 522:25]
    .clock(alu_act_clock),
    .reset(alu_act_reset),
    .io_act_op(alu_act_io_act_op),
    .io_act_en(alu_act_io_act_en),
    .io_i_data_data_0(alu_act_io_i_data_data_0),
    .io_i_data_data_1(alu_act_io_i_data_data_1),
    .io_i_data_data_2(alu_act_io_i_data_data_2),
    .io_i_data_data_3(alu_act_io_i_data_data_3),
    .io_i_data_data_4(alu_act_io_i_data_data_4),
    .io_i_data_data_5(alu_act_io_i_data_data_5),
    .io_i_data_data_6(alu_act_io_i_data_data_6),
    .io_i_data_data_7(alu_act_io_i_data_data_7),
    .io_o_data_data_0(alu_act_io_o_data_data_0),
    .io_o_data_data_1(alu_act_io_o_data_data_1),
    .io_o_data_data_2(alu_act_io_o_data_data_2),
    .io_o_data_data_3(alu_act_io_o_data_data_3),
    .io_o_data_data_4(alu_act_io_o_data_data_4),
    .io_o_data_data_5(alu_act_io_o_data_data_5),
    .io_o_data_data_6(alu_act_io_o_data_data_6),
    .io_o_data_data_7(alu_act_io_o_data_data_7)
  );
  assign io_resize_load = control_io_resize_load; // @[Accel_all.scala 237:19]
  assign io_yolo_finish = control_io_yolo_finish; // @[Accel_all.scala 236:19]
  assign io_conv_finish = control_io_conv_finish; // @[Accel_all.scala 189:40 223:29]
  assign io_dma_raddr = dma_ddr2accel_io_dma_raddr; // @[Accel_all.scala 296:18]
  assign io_dma_rareq = dma_ddr2accel_io_dma_rareq; // @[Accel_all.scala 295:18]
  assign io_dma_rsize = dma_ddr2accel_io_dma_rsize; // @[Accel_all.scala 297:18]
  assign io_dma_rready = 1'h1; // @[Accel_all.scala 294:19]
  assign io_dma_waddr = dma_accel2ddr_io_dma_waddr; // @[Accel_all.scala 278:18]
  assign io_dma_wareq = dma_accel2ddr_io_dma_wareq; // @[Accel_all.scala 275:18]
  assign io_dma_wsize = dma_accel2ddr_io_dma_wsize; // @[Accel_all.scala 279:18]
  assign io_dma_wdata = dma_accel2ddr_io_dma_wdata; // @[Accel_all.scala 280:18]
  assign io_dma_wvalid = dma_accel2ddr_io_dma_wvalid; // @[Accel_all.scala 273:19]
  assign control_clock = clock;
  assign control_reset = reset;
  assign control_io_ap_done = generate_ctrl_signal_io_ap_done; // @[Accel_all.scala 320:13 97:23]
  assign control_io_pool_finish_edge = accel_top_io_pool_finish; // @[Accel_all.scala 215:32 449:21]
  assign control_signal_clock = clock;
  assign control_signal_reset = reset;
  assign control_signal_io_shutdown = generate_ctrl_signal_io_conv_shutdown; // @[Accel_all.scala 317:19 95:29]
  assign control_signal_io_skip_act = reg_0[17]; // @[Accel_all.scala 140:20]
  assign control_signal_io_conv_col = reg_8[9:0]; // @[Accel_all.scala 177:17]
  assign control_signal_io_conv_row = {{2'd0}, row}; // @[Accel_all.scala 246:32]
  assign control_signal_io_s_mod = reg_0[18]; // @[Accel_all.scala 141:17]
  assign control_signal_io_kernal = reg_2[24]; // @[Accel_all.scala 153:21]
  assign control_signal_io_pad_top = pad_cfg[2] & pad_cfg[0]; // @[Accel_all.scala 210:24]
  assign control_signal_io_pad_bottom = pad_cfg[2] & pad_cfg[1]; // @[Accel_all.scala 211:27]
  assign control_signal_io_pad_left_and_right = pad_cfg[2]; // @[Accel_all.scala 212:32]
  assign control_signal_io_pad_size = pad_cfg[2]; // @[Accel_all.scala 213:22]
  assign dma_accel2ddr_clock = clock;
  assign dma_accel2ddr_reset = reset;
  assign dma_accel2ddr_io_send_enable = reg_0[1]; // @[Accel_all.scala 129:25]
  assign dma_accel2ddr_io_dma_addr = control_io_reg6; // @[Accel_all.scala 230:10 50:21]
  assign dma_accel2ddr_io_dma_len = reg_7[18:3]; // @[Accel_all.scala 170:35]
  assign dma_accel2ddr_io_dma_wbusy = io_dma_wbusy; // @[Accel_all.scala 274:32]
  assign dma_accel2ddr_io_dma_wready = io_dma_wready; // @[Accel_all.scala 276:33]
  assign dma_accel2ddr_io_addr_start = {{1'd0}, addr_start}; // @[Accel_all.scala 285:33]
  assign dma_accel2ddr_io_addr_end = {{1'd0}, addr_end}; // @[Accel_all.scala 286:31]
  assign dma_accel2ddr_io_read_data = accel_top_io_ofm_out_bundle; // @[Accel_all.scala 352:28 411:20]
  assign dma_ddr2accel_clock = clock;
  assign dma_ddr2accel_reset = reset;
  assign dma_ddr2accel_io_recv_enable = reg_0[0]; // @[Accel_all.scala 128:25]
  assign dma_ddr2accel_io_dma_addr = control_io_reg4; // @[Accel_all.scala 228:10 48:21]
  assign dma_ddr2accel_io_dma_len = reg_5[18:3]; // @[Accel_all.scala 168:35]
  assign dma_ddr2accel_io_dma_rvalid = io_dma_rvalid; // @[Accel_all.scala 291:33]
  assign dma_ddr2accel_io_dma_rbusy = io_dma_rbusy; // @[Accel_all.scala 292:32]
  assign dma_ddr2accel_io_dma_rdata = io_dma_rdata; // @[Accel_all.scala 293:32]
  assign generate_ctrl_signal_clock = clock;
  assign generate_ctrl_signal_reset = reset;
  assign generate_ctrl_signal_io_recv_enable = reg_0[0]; // @[Accel_all.scala 128:25]
  assign generate_ctrl_signal_io_send_enable = reg_0[1]; // @[Accel_all.scala 129:25]
  assign generate_ctrl_signal_io_conv_start = reg_0[4]; // @[Accel_all.scala 131:24]
  assign generate_ctrl_signal_io_bottleneck_add_enable = reg_0[19]; // @[Accel_all.scala 142:33]
  assign generate_ctrl_signal_io_recv_done = dma_ddr2accel_io_recv_done; // @[Accel_all.scala 299:15 69:25]
  assign generate_ctrl_signal_io_send_done = dma_accel2ddr_io_send_done; // @[Accel_all.scala 282:15 59:25]
  assign generate_ctrl_signal_io_conv_done = yolo_cls_en ? yolo_cls_finish : ofm_done; // @[Accel_all.scala 115:21]
  assign generate_ctrl_signal_io_bottleneck_add_done = accel_top_io_bottleneck_add_finish; // @[Accel_all.scala 216:36 450:26]
  assign generate_ctrl_signal_io_task_valid = reg_0[9]; // @[Accel_all.scala 136:24]
  assign axis_buf_sel_m_io_axis_buf_sel = reg_0[3:2]; // @[Accel_all.scala 130:26]
  assign axis_buf_sel_m_io_write_data = dma_ddr2accel_io_write_data; // @[Accel_all.scala 303:16 73:26]
  assign axis_buf_sel_m_io_write_enable = dma_ddr2accel_io_write_enable; // @[Accel_all.scala 304:18 74:28]
  assign accel_top_clock = clock;
  assign accel_top_reset = reset;
  assign accel_top_io_sel = reg_0[12:10]; // @[Accel_all.scala 137:21]
  assign accel_top_io_ifmbuf_bram_addr_read_s1 = control_signal_io_ifmbuf_bram_addr_read_s1; // @[Accel_all.scala 102:40 250:29]
  assign accel_top_io_ifmbuf_bram_addr_read_sel_s1 = control_signal_io_ifmbuf_addr_read_sel_s1; // @[Accel_all.scala 103:39 251:28]
  assign accel_top_io_ifmbuf_bram_addr_read_s2_singal = control_signal_io_ifmbuf_bram_addr_read_s2_singal; // @[Accel_all.scala 104:47 252:36]
  assign accel_top_io_ifmbuf_bram_addr_read_s2_double = control_signal_io_ifmbuf_bram_addr_read_s2_double; // @[Accel_all.scala 105:47 253:36]
  assign accel_top_io_ifmbuf_sel = reg_0[8]; // @[Accel_all.scala 135:24]
  assign accel_top_io_ifmbuf_bram_en_write = axis_buf_sel_m_io_write_enable_ifm; // @[Accel_all.scala 329:22 80:32]
  assign accel_top_io_recv_done = dma_ddr2accel_io_recv_done; // @[Accel_all.scala 299:15 69:25]
  assign accel_top_io_weightbuf_waddr_clear = ~weightbuf_waddr_clear_REG & task_valid; // @[utils.scala 10:27]
  assign accel_top_io_weightbuf_bram_en_write = axis_buf_sel_m_io_write_enable_weight; // @[Accel_all.scala 332:25 83:35]
  assign accel_top_io_weightbuf_read_addr = reg_3[6:0]; // @[Accel_all.scala 157:36]
  assign accel_top_io_kernal = reg_2[24]; // @[Accel_all.scala 153:21]
  assign accel_top_io_weight_sel = reg_3[15:13]; // @[Accel_all.scala 159:25]
  assign accel_top_io_biasbuf_waddr_clear = ~biasbuf_waddr_clear_REG & task_valid; // @[utils.scala 10:27]
  assign accel_top_io_biasbuf_bram_en_write = axis_buf_sel_m_io_write_enable_bias; // @[Accel_all.scala 335:23 86:33]
  assign accel_top_io_biasbuf_read_addr = reg_3[22:16]; // @[Accel_all.scala 158:34]
  assign accel_top_io_acc_read_en = control_signal_io_acc_read_en; // @[Accel_all.scala 108:27 256:16]
  assign accel_top_io_acc_write_en = control_signal_io_acc_write_en; // @[Accel_all.scala 109:28 257:17]
  assign accel_top_io_acc_read_addr = control_signal_io_acc_read_addr; // @[Accel_all.scala 106:29 254:18]
  assign accel_top_io_acc_write_addr = control_signal_io_acc_write_addr; // @[Accel_all.scala 107:30 255:19]
  assign accel_top_io_acc_prev_data_zero = reg_0[6]; // @[Accel_all.scala 133:24]
  assign accel_top_io_acc_curr_data_zero = control_signal_io_acc_curr_data_zero; // @[Accel_all.scala 110:34 258:23]
  assign accel_top_io_ofmbuf_bram_en_write = yolo_cls_en ? yolo_ofm_write_en_after : ofm_valid; // @[Accel_all.scala 408:45]
  assign accel_top_io_ofmbuf_bram_write_addr = _accel_top_io_ofmbuf_bram_write_addr_T[11:0]; // @[Accel_all.scala 409:41]
  assign accel_top_io_ofmbuf_bram_read_addr = {{52'd0}, _accel_top_io_ofmbuf_bram_read_addr_T}; // @[Accel_all.scala 410:40]
  assign accel_top_io_col = reg_8[9:0]; // @[Accel_all.scala 177:17]
  assign accel_top_io_row = {{2'd0}, row}; // @[Accel_all.scala 436:22]
  assign accel_top_io_pad_top = pad_cfg[2] & pad_cfg[0]; // @[Accel_all.scala 210:24]
  assign accel_top_io_pad_bottom = pad_cfg[2] & pad_cfg[1]; // @[Accel_all.scala 211:27]
  assign accel_top_io_pad_left_and_right = pad_cfg[2]; // @[Accel_all.scala 212:32]
  assign accel_top_io_zero_pad_valid_s2 = control_signal_io_zero_pad_valid_s2; // @[Accel_all.scala 209:31 267:23]
  assign accel_top_io_zero_pad_valid_s1 = control_signal_io_zero_pad_valid_s1; // @[Accel_all.scala 208:33 268:23]
  assign accel_top_io_scale = reg_1[15:0]; // @[Accel_all.scala 146:20]
  assign accel_top_io_shift = reg_1[19:16]; // @[Accel_all.scala 147:20]
  assign accel_top_io_zero_point_in = reg_2[7:0]; // @[Accel_all.scala 150:30]
  assign accel_top_io_zero_point_out = reg_2[15:8]; // @[Accel_all.scala 151:31]
  assign accel_top_io_zero_point_A_act = reg_2[23:16]; // @[Accel_all.scala 152:31]
  assign accel_top_io_ifm_in_0 = write_data_ifm[7:0]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_1 = write_data_ifm[15:8]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_2 = write_data_ifm[23:16]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_3 = write_data_ifm[31:24]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_4 = write_data_ifm[39:32]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_5 = write_data_ifm[47:40]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_6 = write_data_ifm[55:48]; // @[Accel_all.scala 342:34]
  assign accel_top_io_ifm_in_7 = write_data_ifm[63:56]; // @[Accel_all.scala 342:34]
  assign accel_top_io_weight_in_0 = write_data_weight[7:0]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_1 = write_data_weight[15:8]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_2 = write_data_weight[23:16]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_3 = write_data_weight[31:24]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_4 = write_data_weight[39:32]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_5 = write_data_weight[47:40]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_6 = write_data_weight[55:48]; // @[Accel_all.scala 346:40]
  assign accel_top_io_weight_in_7 = write_data_weight[63:56]; // @[Accel_all.scala 346:40]
  assign accel_top_io_bias_in = write_data_bias[17:0]; // @[Accel_all.scala 348:21 349:12]
  assign accel_top_io_bias_valid = reg_0[7]; // @[Accel_all.scala 134:23]
  assign accel_top_io_skip_act = reg_0[17]; // @[Accel_all.scala 140:20]
  assign accel_top_io_pool_enable = reg_0[5]; // @[Accel_all.scala 132:25]
  assign accel_top_io_upsample_enable = reg_0[16]; // @[Accel_all.scala 139:29]
  assign accel_top_io_bottleneck_add_enable = reg_0[19]; // @[Accel_all.scala 142:33]
  assign accel_top_io_s_mod = reg_0[18]; // @[Accel_all.scala 141:17]
  assign accel_top_io_act_outdata_0 = quant_io_o_data_0; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_1 = quant_io_o_data_1; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_2 = quant_io_o_data_2; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_3 = quant_io_o_data_3; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_4 = quant_io_o_data_4; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_5 = quant_io_o_data_5; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_6 = quant_io_o_data_6; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_act_outdata_7 = quant_io_o_data_7; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_0 = quant_io_o_data_0; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_1 = quant_io_o_data_1; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_2 = quant_io_o_data_2; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_3 = quant_io_o_data_3; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_4 = quant_io_o_data_4; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_5 = quant_io_o_data_5; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_6 = quant_io_o_data_6; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_bn_add_result_7 = quant_io_o_data_7; // @[Accel_all.scala 362:25 517:15]
  assign accel_top_io_yolo_cls_en = reg_8[16]; // @[Accel_all.scala 179:25]
  assign accel_top_io_yolo_cls_data_after_compare = yolo_io_ofm_write_data_after; // @[Accel_all.scala 371:41 474:33]
  assign yolo_clock = clock;
  assign yolo_reset = reset;
  assign yolo_io_yolo_layer_cls_en = reg_8[16]; // @[Accel_all.scala 179:25]
  assign yolo_io_yolo_current_cls_detect_layer = reg_8[19:18]; // @[Accel_all.scala 181:46]
  assign yolo_io_yolo_layer_cls_div_cnt = reg_8[23:20]; // @[Accel_all.scala 182:39]
  assign yolo_io_ofm_write_data_before = accel_top_io_yolo_cls_data_before_compare; // @[Accel_all.scala 370:42 457:34]
  assign yolo_io_ofm_write_en_before = ofm_valid & ~ofm_write_disable; // @[Accel_all.scala 473:46]
  assign yolo_io_data_after_sigmoid = alu_act_out_0[23:0]; // @[Accel_all.scala 481:46]
  assign dequant_clock = clock;
  assign dequant_reset = reset;
  assign dequant_io_en = _act_op_T | bn_add_working; // @[Accel_all.scala 495:31]
  assign dequant_io_i_data_0 = _act_op_T ? act_indata_0 : _dequant_in_0_T_4; // @[Mux.scala 101:16]
  assign dequant_io_i_data_1 = _act_op_T ? act_indata_1 : _dequant_in_1_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_2 = _act_op_T ? act_indata_2 : _dequant_in_2_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_3 = _act_op_T ? act_indata_3 : _dequant_in_3_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_4 = _act_op_T ? act_indata_4 : _dequant_in_4_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_5 = _act_op_T ? act_indata_5 : _dequant_in_5_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_6 = _act_op_T ? act_indata_6 : _dequant_in_6_T_2; // @[Mux.scala 101:16]
  assign dequant_io_i_data_7 = _act_op_T ? act_indata_7 : _dequant_in_7_T_2; // @[Mux.scala 101:16]
  assign dequant_io_scale = control_io_reg9; // @[Accel_all.scala 233:10 54:21]
  assign dequant_io_zero_point = reg_2[15:8]; // @[Accel_all.scala 151:31]
  assign dequant_extra_clock = clock;
  assign dequant_extra_reset = reset;
  assign dequant_extra_io_en = _act_op_T | bn_add_working; // @[Accel_all.scala 502:37]
  assign dequant_extra_io_i_data_0 = accel_top_io_bn_add_in1_0; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_1 = accel_top_io_bn_add_in1_1; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_2 = accel_top_io_bn_add_in1_2; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_3 = accel_top_io_bn_add_in1_3; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_4 = accel_top_io_bn_add_in1_4; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_5 = accel_top_io_bn_add_in1_5; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_6 = accel_top_io_bn_add_in1_6; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_i_data_7 = accel_top_io_bn_add_in1_7; // @[Accel_all.scala 359:26 453:16]
  assign dequant_extra_io_scale = dequant_extra_scala; // @[Accel_all.scala 505:28]
  assign dequant_extra_io_zero_point = dequant_extra_zero_point; // @[Accel_all.scala 506:33]
  assign bn_add_float_result_0_adder_clock = clock;
  assign bn_add_float_result_0_adder_reset = reset;
  assign bn_add_float_result_0_adder_io_x = dequant_io_o_data_0; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_0_adder_io_y = dequant_extra_io_o_data_0; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_0_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_1_adder_clock = clock;
  assign bn_add_float_result_1_adder_reset = reset;
  assign bn_add_float_result_1_adder_io_x = dequant_io_o_data_1; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_1_adder_io_y = dequant_extra_io_o_data_1; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_1_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_2_adder_clock = clock;
  assign bn_add_float_result_2_adder_reset = reset;
  assign bn_add_float_result_2_adder_io_x = dequant_io_o_data_2; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_2_adder_io_y = dequant_extra_io_o_data_2; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_2_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_3_adder_clock = clock;
  assign bn_add_float_result_3_adder_reset = reset;
  assign bn_add_float_result_3_adder_io_x = dequant_io_o_data_3; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_3_adder_io_y = dequant_extra_io_o_data_3; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_3_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_4_adder_clock = clock;
  assign bn_add_float_result_4_adder_reset = reset;
  assign bn_add_float_result_4_adder_io_x = dequant_io_o_data_4; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_4_adder_io_y = dequant_extra_io_o_data_4; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_4_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_5_adder_clock = clock;
  assign bn_add_float_result_5_adder_reset = reset;
  assign bn_add_float_result_5_adder_io_x = dequant_io_o_data_5; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_5_adder_io_y = dequant_extra_io_o_data_5; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_5_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_6_adder_clock = clock;
  assign bn_add_float_result_6_adder_reset = reset;
  assign bn_add_float_result_6_adder_io_x = dequant_io_o_data_6; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_6_adder_io_y = dequant_extra_io_o_data_6; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_6_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign bn_add_float_result_7_adder_clock = clock;
  assign bn_add_float_result_7_adder_reset = reset;
  assign bn_add_float_result_7_adder_io_x = dequant_io_o_data_7; // @[Accel_all.scala 492:34 497:23]
  assign bn_add_float_result_7_adder_io_y = dequant_extra_io_o_data_7; // @[Accel_all.scala 493:45 504:34]
  assign bn_add_float_result_7_adder_io_valid_in = generate_ctrl_signal_io_bn_add_working; // @[Accel_all.scala 217:30 318:20]
  assign quant_clock = clock;
  assign quant_reset = reset;
  assign quant_io_en = _act_op_T | bn_add_working; // @[Accel_all.scala 515:32]
  assign quant_io_i_data_0 = bn_add_working ? bn_add_float_result_0_result_2_bits : alu_act_out_0; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_1 = bn_add_working ? bn_add_float_result_1_result_2_bits : alu_act_out_1; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_2 = bn_add_working ? bn_add_float_result_2_result_2_bits : alu_act_out_2; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_3 = bn_add_working ? bn_add_float_result_3_result_2_bits : alu_act_out_3; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_4 = bn_add_working ? bn_add_float_result_4_result_2_bits : alu_act_out_4; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_5 = bn_add_working ? bn_add_float_result_5_result_2_bits : alu_act_out_5; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_6 = bn_add_working ? bn_add_float_result_6_result_2_bits : alu_act_out_6; // @[Accel_all.scala 516:27]
  assign quant_io_i_data_7 = bn_add_working ? bn_add_float_result_7_result_2_bits : alu_act_out_7; // @[Accel_all.scala 516:27]
  assign quant_io_scale = control_io_reg10; // @[Accel_all.scala 234:11 55:22]
  assign quant_io_zero_point = reg_2[23:16]; // @[Accel_all.scala 152:31]
  assign alu_act_clock = clock;
  assign alu_act_reset = reset;
  assign alu_act_io_act_op = sigmoid_en ? 2'h2 : {{1'd0}, _act_op_T}; // @[Accel_all.scala 463:21]
  assign alu_act_io_act_en = _act_op_T | sigmoid_en; // @[Accel_all.scala 526:38]
  assign alu_act_io_i_data_data_0 = dequant_io_o_data_0; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_1 = dequant_io_o_data_1; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_2 = dequant_io_o_data_2; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_3 = dequant_io_o_data_3; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_4 = dequant_io_o_data_4; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_5 = dequant_io_o_data_5; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_6 = dequant_io_o_data_6; // @[Accel_all.scala 492:34 497:23]
  assign alu_act_io_i_data_data_7 = dequant_io_o_data_7; // @[Accel_all.scala 492:34 497:23]
  always @(posedge clock) begin
    if (reset) begin // @[utils.scala 10:17]
      weightbuf_waddr_clear_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      weightbuf_waddr_clear_REG <= task_valid; // @[utils.scala 10:17]
    end
    if (reset) begin // @[utils.scala 10:17]
      biasbuf_waddr_clear_REG <= 1'h0; // @[utils.scala 10:17]
    end else begin
      biasbuf_waddr_clear_REG <= task_valid; // @[utils.scala 10:17]
    end
    if (reset) begin // @[Reg.scala 35:20]
      dequant_extra_scala_temp <= 32'h0; // @[Reg.scala 35:20]
    end else if (conv_finish_from_control) begin // @[Reg.scala 36:18]
      dequant_extra_scala_temp <= dequant_scala; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      dequant_extra_scala <= 32'h0; // @[Reg.scala 35:20]
    end else if (conv_finish_from_control) begin // @[Reg.scala 36:18]
      dequant_extra_scala <= dequant_extra_scala_temp; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      dequant_extra_zero_point_temp <= 8'h0; // @[Reg.scala 35:20]
    end else if (conv_finish_from_control) begin // @[Reg.scala 36:18]
      dequant_extra_zero_point_temp <= dequant_zero_point; // @[Reg.scala 36:22]
    end
    if (reset) begin // @[Reg.scala 35:20]
      dequant_extra_zero_point <= 8'h0; // @[Reg.scala 35:20]
    end else if (conv_finish_from_control) begin // @[Reg.scala 36:18]
      dequant_extra_zero_point <= dequant_extra_zero_point_temp; // @[Reg.scala 36:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  weightbuf_waddr_clear_REG = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  biasbuf_waddr_clear_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dequant_extra_scala_temp = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dequant_extra_scala = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dequant_extra_zero_point_temp = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  dequant_extra_zero_point = _RAND_5[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
